`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   10:36:36 12/13/2016
// Design Name:   MFCC
// Module Name:   C:/Users/tslab-802-2/Desktop/newtest/FPGA_project - backup1/MFC_REC/simtest.v
// Project Name:  MFC_REC
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: MFCC
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module simtest;

	// Inputs
	reg clk;
	reg [15:0] x_i;
	reg write;
	reg 	  reset;
	reg [16:0] index2=0;
	reg [16:0] index=0;
	// Outputs
	wire [31:0] x_o;
	wire [4:0] out_index;
	wire dv;
	wire vad;
//	wire [3:0] process=0;

	// Instantiate the Unit Under Test (UUT)
	MFCC MFCC(.clk(clk),
	     .sclk(clk),
	     .x_i(x_i), 
	     .write(write),
	     .dv_out(dv), 
	     .out_index(out_index), 
	     .x_o(x_o),
		  .vad(vad));
	
	wire signed [21:0] dnn_out;
	wire dnn_dv;
//	wire signed [16:0]indataA1 = 0;	//16bit
//	wire signed [14:0]indataB1 = 0;	//14bit
	DNN_0117 nnmain (
		 .clk(clk), 
		 .reset(reset), 
		 .vec_in(x_o), 
		 .dv_in(dv), 
		 .vec_out(dnn_out), 
		 .dv_out(dnn_dv)
		 );
		 
		 
	always begin 
		#5
		clk <= ~clk;
		case (index)
default:begin
end
0:begin
x_i <= 19;
end
1:begin
x_i <= 27;
end
2:begin
x_i <= 31;
end
3:begin
x_i <= 72;
end
4:begin
x_i <= 40;
end
5:begin
x_i <= 70;
end
6:begin
x_i <= 24;
end
7:begin
x_i <= 27;
end
8:begin
x_i <= 37;
end
9:begin
x_i <= 30;
end
10:begin
x_i <= 43;
end
11:begin
x_i <= 19;
end
12:begin
x_i <= 19;
end
13:begin
x_i <= 13;
end
14:begin
x_i <= 65524;
end
15:begin
x_i <= 65499;
end
16:begin
x_i <= 65526;
end
17:begin
x_i <= 65515;
end
18:begin
x_i <= 65502;
end
19:begin
x_i <= 65507;
end
20:begin
x_i <= 65490;
end
21:begin
x_i <= 65498;
end
22:begin
x_i <= 65510;
end
23:begin
x_i <= 65482;
end
24:begin
x_i <= 65514;
end
25:begin
x_i <= 65494;
end
26:begin
x_i <= 65466;
end
27:begin
x_i <= 65494;
end
28:begin
x_i <= 65506;
end
29:begin
x_i <= 65521;
end
30:begin
x_i <= 65467;
end
31:begin
x_i <= 65478;
end
32:begin
x_i <= 65498;
end
33:begin
x_i <= 65522;
end
34:begin
x_i <= 65514;
end
35:begin
x_i <= 65516;
end
36:begin
x_i <= 65514;
end
37:begin
x_i <= 65503;
end
38:begin
x_i <= 65533;
end
39:begin
x_i <= 65497;
end
40:begin
x_i <= 65511;
end
41:begin
x_i <= 65490;
end
42:begin
x_i <= 65464;
end
43:begin
x_i <= 65451;
end
44:begin
x_i <= 65473;
end
45:begin
x_i <= 65470;
end
46:begin
x_i <= 65469;
end
47:begin
x_i <= 65482;
end
48:begin
x_i <= 65450;
end
49:begin
x_i <= 65457;
end
50:begin
x_i <= 65434;
end
51:begin
x_i <= 65451;
end
52:begin
x_i <= 65462;
end
53:begin
x_i <= 65424;
end
54:begin
x_i <= 65413;
end
55:begin
x_i <= 65452;
end
56:begin
x_i <= 65460;
end
57:begin
x_i <= 65454;
end
58:begin
x_i <= 65434;
end
59:begin
x_i <= 65474;
end
60:begin
x_i <= 65473;
end
61:begin
x_i <= 65449;
end
62:begin
x_i <= 65485;
end
63:begin
x_i <= 65443;
end
64:begin
x_i <= 65451;
end
65:begin
x_i <= 65470;
end
66:begin
x_i <= 65486;
end
67:begin
x_i <= 65474;
end
68:begin
x_i <= 65489;
end
69:begin
x_i <= 65482;
end
70:begin
x_i <= 65471;
end
71:begin
x_i <= 65494;
end
72:begin
x_i <= 65478;
end
73:begin
x_i <= 65501;
end
74:begin
x_i <= 65521;
end
75:begin
x_i <= 5;
end
76:begin
x_i <= 37;
end
77:begin
x_i <= 62;
end
78:begin
x_i <= 68;
end
79:begin
x_i <= 70;
end
80:begin
x_i <= 51;
end
81:begin
x_i <= 65535;
end
82:begin
x_i <= 5;
end
83:begin
x_i <= 33;
end
84:begin
x_i <= 2;
end
85:begin
x_i <= 95;
end
86:begin
x_i <= 82;
end
87:begin
x_i <= 86;
end
88:begin
x_i <= 147;
end
89:begin
x_i <= 137;
end
90:begin
x_i <= 124;
end
91:begin
x_i <= 78;
end
92:begin
x_i <= 35;
end
93:begin
x_i <= 56;
end
94:begin
x_i <= 16;
end
95:begin
x_i <= 65481;
end
96:begin
x_i <= 65466;
end
97:begin
x_i <= 65420;
end
98:begin
x_i <= 65421;
end
99:begin
x_i <= 65444;
end
100:begin
x_i <= 65471;
end
101:begin
x_i <= 65520;
end
102:begin
x_i <= 65530;
end
103:begin
x_i <= 33;
end
104:begin
x_i <= 37;
end
105:begin
x_i <= 32;
end
106:begin
x_i <= 30;
end
107:begin
x_i <= 17;
end
108:begin
x_i <= 65526;
end
109:begin
x_i <= 65482;
end
110:begin
x_i <= 65456;
end
111:begin
x_i <= 65531;
end
112:begin
x_i <= 65505;
end
113:begin
x_i <= 65514;
end
114:begin
x_i <= 65523;
end
115:begin
x_i <= 65516;
end
116:begin
x_i <= 65530;
end
117:begin
x_i <= 65521;
end
118:begin
x_i <= 65496;
end
119:begin
x_i <= 65487;
end
120:begin
x_i <= 65469;
end
121:begin
x_i <= 65488;
end
122:begin
x_i <= 65500;
end
123:begin
x_i <= 65508;
end
124:begin
x_i <= 65485;
end
125:begin
x_i <= 65479;
end
126:begin
x_i <= 65461;
end
127:begin
x_i <= 65453;
end
128:begin
x_i <= 65436;
end
129:begin
x_i <= 65399;
end
130:begin
x_i <= 65427;
end
131:begin
x_i <= 65424;
end
132:begin
x_i <= 65437;
end
133:begin
x_i <= 65476;
end
134:begin
x_i <= 65517;
end
135:begin
x_i <= 65529;
end
136:begin
x_i <= 65516;
end
137:begin
x_i <= 65495;
end
138:begin
x_i <= 65434;
end
139:begin
x_i <= 65386;
end
140:begin
x_i <= 65387;
end
141:begin
x_i <= 65374;
end
142:begin
x_i <= 65414;
end
143:begin
x_i <= 65430;
end
144:begin
x_i <= 65467;
end
145:begin
x_i <= 65489;
end
146:begin
x_i <= 65502;
end
147:begin
x_i <= 65520;
end
148:begin
x_i <= 65485;
end
149:begin
x_i <= 65458;
end
150:begin
x_i <= 65437;
end
151:begin
x_i <= 65440;
end
152:begin
x_i <= 65473;
end
153:begin
x_i <= 65500;
end
154:begin
x_i <= 65532;
end
155:begin
x_i <= 54;
end
156:begin
x_i <= 82;
end
157:begin
x_i <= 85;
end
158:begin
x_i <= 102;
end
159:begin
x_i <= 87;
end
160:begin
x_i <= 24;
end
161:begin
x_i <= 69;
end
162:begin
x_i <= 48;
end
163:begin
x_i <= 50;
end
164:begin
x_i <= 95;
end
165:begin
x_i <= 113;
end
166:begin
x_i <= 138;
end
167:begin
x_i <= 186;
end
168:begin
x_i <= 217;
end
169:begin
x_i <= 167;
end
170:begin
x_i <= 128;
end
171:begin
x_i <= 110;
end
172:begin
x_i <= 38;
end
173:begin
x_i <= 65524;
end
174:begin
x_i <= 65429;
end
175:begin
x_i <= 65345;
end
176:begin
x_i <= 65336;
end
177:begin
x_i <= 65366;
end
178:begin
x_i <= 65468;
end
179:begin
x_i <= 65526;
end
180:begin
x_i <= 51;
end
181:begin
x_i <= 73;
end
182:begin
x_i <= 98;
end
183:begin
x_i <= 58;
end
184:begin
x_i <= 13;
end
185:begin
x_i <= 65527;
end
186:begin
x_i <= 65474;
end
187:begin
x_i <= 65411;
end
188:begin
x_i <= 65378;
end
189:begin
x_i <= 65439;
end
190:begin
x_i <= 65527;
end
191:begin
x_i <= 65526;
end
192:begin
x_i <= 65514;
end
193:begin
x_i <= 43;
end
194:begin
x_i <= 16;
end
195:begin
x_i <= 65481;
end
196:begin
x_i <= 65464;
end
197:begin
x_i <= 65463;
end
198:begin
x_i <= 65457;
end
199:begin
x_i <= 65435;
end
200:begin
x_i <= 65454;
end
201:begin
x_i <= 65499;
end
202:begin
x_i <= 25;
end
203:begin
x_i <= 65534;
end
204:begin
x_i <= 65500;
end
205:begin
x_i <= 65478;
end
206:begin
x_i <= 65452;
end
207:begin
x_i <= 65378;
end
208:begin
x_i <= 65376;
end
209:begin
x_i <= 65401;
end
210:begin
x_i <= 65403;
end
211:begin
x_i <= 65448;
end
212:begin
x_i <= 1;
end
213:begin
x_i <= 66;
end
214:begin
x_i <= 59;
end
215:begin
x_i <= 24;
end
216:begin
x_i <= 65483;
end
217:begin
x_i <= 65419;
end
218:begin
x_i <= 65359;
end
219:begin
x_i <= 65330;
end
220:begin
x_i <= 65371;
end
221:begin
x_i <= 65376;
end
222:begin
x_i <= 65428;
end
223:begin
x_i <= 65468;
end
224:begin
x_i <= 65500;
end
225:begin
x_i <= 65520;
end
226:begin
x_i <= 65508;
end
227:begin
x_i <= 65479;
end
228:begin
x_i <= 65468;
end
229:begin
x_i <= 65441;
end
230:begin
x_i <= 65446;
end
231:begin
x_i <= 65470;
end
232:begin
x_i <= 65495;
end
233:begin
x_i <= 15;
end
234:begin
x_i <= 63;
end
235:begin
x_i <= 83;
end
236:begin
x_i <= 101;
end
237:begin
x_i <= 68;
end
238:begin
x_i <= 40;
end
239:begin
x_i <= 30;
end
240:begin
x_i <= 36;
end
241:begin
x_i <= 64;
end
242:begin
x_i <= 62;
end
243:begin
x_i <= 110;
end
244:begin
x_i <= 157;
end
245:begin
x_i <= 199;
end
246:begin
x_i <= 216;
end
247:begin
x_i <= 242;
end
248:begin
x_i <= 184;
end
249:begin
x_i <= 213;
end
250:begin
x_i <= 132;
end
251:begin
x_i <= 58;
end
252:begin
x_i <= 65522;
end
253:begin
x_i <= 65346;
end
254:begin
x_i <= 65175;
end
255:begin
x_i <= 65166;
end
256:begin
x_i <= 65259;
end
257:begin
x_i <= 65440;
end
258:begin
x_i <= 17;
end
259:begin
x_i <= 72;
end
260:begin
x_i <= 195;
end
261:begin
x_i <= 202;
end
262:begin
x_i <= 106;
end
263:begin
x_i <= 44;
end
264:begin
x_i <= 65505;
end
265:begin
x_i <= 65380;
end
266:begin
x_i <= 65293;
end
267:begin
x_i <= 65302;
end
268:begin
x_i <= 65396;
end
269:begin
x_i <= 65515;
end
270:begin
x_i <= 65533;
end
271:begin
x_i <= 50;
end
272:begin
x_i <= 94;
end
273:begin
x_i <= 39;
end
274:begin
x_i <= 65509;
end
275:begin
x_i <= 65429;
end
276:begin
x_i <= 65427;
end
277:begin
x_i <= 65393;
end
278:begin
x_i <= 65399;
end
279:begin
x_i <= 65496;
end
280:begin
x_i <= 65535;
end
281:begin
x_i <= 33;
end
282:begin
x_i <= 18;
end
283:begin
x_i <= 9;
end
284:begin
x_i <= 65483;
end
285:begin
x_i <= 65392;
end
286:begin
x_i <= 65324;
end
287:begin
x_i <= 65314;
end
288:begin
x_i <= 65331;
end
289:begin
x_i <= 65407;
end
290:begin
x_i <= 65519;
end
291:begin
x_i <= 99;
end
292:begin
x_i <= 120;
end
293:begin
x_i <= 88;
end
294:begin
x_i <= 52;
end
295:begin
x_i <= 65476;
end
296:begin
x_i <= 65346;
end
297:begin
x_i <= 65268;
end
298:begin
x_i <= 65257;
end
299:begin
x_i <= 65232;
end
300:begin
x_i <= 65338;
end
301:begin
x_i <= 65436;
end
302:begin
x_i <= 65526;
end
303:begin
x_i <= 31;
end
304:begin
x_i <= 27;
end
305:begin
x_i <= 13;
end
306:begin
x_i <= 65492;
end
307:begin
x_i <= 65440;
end
308:begin
x_i <= 65449;
end
309:begin
x_i <= 65460;
end
310:begin
x_i <= 65458;
end
311:begin
x_i <= 65505;
end
312:begin
x_i <= 65532;
end
313:begin
x_i <= 23;
end
314:begin
x_i <= 77;
end
315:begin
x_i <= 81;
end
316:begin
x_i <= 58;
end
317:begin
x_i <= 66;
end
318:begin
x_i <= 45;
end
319:begin
x_i <= 51;
end
320:begin
x_i <= 95;
end
321:begin
x_i <= 80;
end
322:begin
x_i <= 190;
end
323:begin
x_i <= 197;
end
324:begin
x_i <= 232;
end
325:begin
x_i <= 274;
end
326:begin
x_i <= 255;
end
327:begin
x_i <= 246;
end
328:begin
x_i <= 250;
end
329:begin
x_i <= 201;
end
330:begin
x_i <= 161;
end
331:begin
x_i <= 4;
end
332:begin
x_i <= 65312;
end
333:begin
x_i <= 65107;
end
334:begin
x_i <= 65016;
end
335:begin
x_i <= 65170;
end
336:begin
x_i <= 65459;
end
337:begin
x_i <= 56;
end
338:begin
x_i <= 157;
end
339:begin
x_i <= 251;
end
340:begin
x_i <= 337;
end
341:begin
x_i <= 217;
end
342:begin
x_i <= 82;
end
343:begin
x_i <= 65439;
end
344:begin
x_i <= 65300;
end
345:begin
x_i <= 65176;
end
346:begin
x_i <= 65155;
end
347:begin
x_i <= 65332;
end
348:begin
x_i <= 65488;
end
349:begin
x_i <= 54;
end
350:begin
x_i <= 110;
end
351:begin
x_i <= 148;
end
352:begin
x_i <= 134;
end
353:begin
x_i <= 48;
end
354:begin
x_i <= 65425;
end
355:begin
x_i <= 65366;
end
356:begin
x_i <= 65343;
end
357:begin
x_i <= 65388;
end
358:begin
x_i <= 65396;
end
359:begin
x_i <= 14;
end
360:begin
x_i <= 82;
end
361:begin
x_i <= 55;
end
362:begin
x_i <= 5;
end
363:begin
x_i <= 65467;
end
364:begin
x_i <= 65365;
end
365:begin
x_i <= 65273;
end
366:begin
x_i <= 65249;
end
367:begin
x_i <= 65325;
end
368:begin
x_i <= 65434;
end
369:begin
x_i <= 13;
end
370:begin
x_i <= 123;
end
371:begin
x_i <= 191;
end
372:begin
x_i <= 129;
end
373:begin
x_i <= 40;
end
374:begin
x_i <= 65419;
end
375:begin
x_i <= 65332;
end
376:begin
x_i <= 65225;
end
377:begin
x_i <= 65207;
end
378:begin
x_i <= 65240;
end
379:begin
x_i <= 65346;
end
380:begin
x_i <= 65457;
end
381:begin
x_i <= 65495;
end
382:begin
x_i <= 10;
end
383:begin
x_i <= 22;
end
384:begin
x_i <= 1;
end
385:begin
x_i <= 65481;
end
386:begin
x_i <= 65468;
end
387:begin
x_i <= 65482;
end
388:begin
x_i <= 65454;
end
389:begin
x_i <= 65474;
end
390:begin
x_i <= 65508;
end
391:begin
x_i <= 65517;
end
392:begin
x_i <= 65521;
end
393:begin
x_i <= 25;
end
394:begin
x_i <= 31;
end
395:begin
x_i <= 46;
end
396:begin
x_i <= 59;
end
397:begin
x_i <= 87;
end
398:begin
x_i <= 126;
end
399:begin
x_i <= 143;
end
400:begin
x_i <= 152;
end
401:begin
x_i <= 217;
end
402:begin
x_i <= 264;
end
403:begin
x_i <= 270;
end
404:begin
x_i <= 297;
end
405:begin
x_i <= 322;
end
406:begin
x_i <= 289;
end
407:begin
x_i <= 323;
end
408:begin
x_i <= 273;
end
409:begin
x_i <= 219;
end
410:begin
x_i <= 75;
end
411:begin
x_i <= 65161;
end
412:begin
x_i <= 64832;
end
413:begin
x_i <= 64940;
end
414:begin
x_i <= 65245;
end
415:begin
x_i <= 5;
end
416:begin
x_i <= 91;
end
417:begin
x_i <= 252;
end
418:begin
x_i <= 490;
end
419:begin
x_i <= 471;
end
420:begin
x_i <= 249;
end
421:begin
x_i <= 51;
end
422:begin
x_i <= 65398;
end
423:begin
x_i <= 65146;
end
424:begin
x_i <= 64974;
end
425:begin
x_i <= 65080;
end
426:begin
x_i <= 65393;
end
427:begin
x_i <= 23;
end
428:begin
x_i <= 111;
end
429:begin
x_i <= 225;
end
430:begin
x_i <= 295;
end
431:begin
x_i <= 184;
end
432:begin
x_i <= 29;
end
433:begin
x_i <= 65393;
end
434:begin
x_i <= 65336;
end
435:begin
x_i <= 65292;
end
436:begin
x_i <= 65327;
end
437:begin
x_i <= 65424;
end
438:begin
x_i <= 51;
end
439:begin
x_i <= 118;
end
440:begin
x_i <= 50;
end
441:begin
x_i <= 65504;
end
442:begin
x_i <= 65459;
end
443:begin
x_i <= 65303;
end
444:begin
x_i <= 65198;
end
445:begin
x_i <= 65257;
end
446:begin
x_i <= 65359;
end
447:begin
x_i <= 65437;
end
448:begin
x_i <= 65526;
end
449:begin
x_i <= 88;
end
450:begin
x_i <= 192;
end
451:begin
x_i <= 112;
end
452:begin
x_i <= 23;
end
453:begin
x_i <= 65465;
end
454:begin
x_i <= 65318;
end
455:begin
x_i <= 65191;
end
456:begin
x_i <= 65142;
end
457:begin
x_i <= 65220;
end
458:begin
x_i <= 65336;
end
459:begin
x_i <= 65359;
end
460:begin
x_i <= 65453;
end
461:begin
x_i <= 88;
end
462:begin
x_i <= 80;
end
463:begin
x_i <= 35;
end
464:begin
x_i <= 11;
end
465:begin
x_i <= 65517;
end
466:begin
x_i <= 65475;
end
467:begin
x_i <= 65457;
end
468:begin
x_i <= 65483;
end
469:begin
x_i <= 16;
end
470:begin
x_i <= 26;
end
471:begin
x_i <= 65524;
end
472:begin
x_i <= 24;
end
473:begin
x_i <= 62;
end
474:begin
x_i <= 40;
end
475:begin
x_i <= 62;
end
476:begin
x_i <= 65;
end
477:begin
x_i <= 128;
end
478:begin
x_i <= 215;
end
479:begin
x_i <= 248;
end
480:begin
x_i <= 310;
end
481:begin
x_i <= 329;
end
482:begin
x_i <= 326;
end
483:begin
x_i <= 336;
end
484:begin
x_i <= 324;
end
485:begin
x_i <= 289;
end
486:begin
x_i <= 277;
end
487:begin
x_i <= 160;
end
488:begin
x_i <= 65258;
end
489:begin
x_i <= 64769;
end
490:begin
x_i <= 64697;
end
491:begin
x_i <= 65063;
end
492:begin
x_i <= 65501;
end
493:begin
x_i <= 67;
end
494:begin
x_i <= 171;
end
495:begin
x_i <= 501;
end
496:begin
x_i <= 603;
end
497:begin
x_i <= 415;
end
498:begin
x_i <= 122;
end
499:begin
x_i <= 65480;
end
500:begin
x_i <= 65209;
end
501:begin
x_i <= 64943;
end
502:begin
x_i <= 64911;
end
503:begin
x_i <= 65196;
end
504:begin
x_i <= 65526;
end
505:begin
x_i <= 92;
end
506:begin
x_i <= 194;
end
507:begin
x_i <= 331;
end
508:begin
x_i <= 332;
end
509:begin
x_i <= 156;
end
510:begin
x_i <= 65458;
end
511:begin
x_i <= 65363;
end
512:begin
x_i <= 65293;
end
513:begin
x_i <= 65241;
end
514:begin
x_i <= 65342;
end
515:begin
x_i <= 65524;
end
516:begin
x_i <= 95;
end
517:begin
x_i <= 68;
end
518:begin
x_i <= 65521;
end
519:begin
x_i <= 65473;
end
520:begin
x_i <= 65340;
end
521:begin
x_i <= 65231;
end
522:begin
x_i <= 65146;
end
523:begin
x_i <= 65191;
end
524:begin
x_i <= 65360;
end
525:begin
x_i <= 65456;
end
526:begin
x_i <= 34;
end
527:begin
x_i <= 174;
end
528:begin
x_i <= 225;
end
529:begin
x_i <= 155;
end
530:begin
x_i <= 23;
end
531:begin
x_i <= 65421;
end
532:begin
x_i <= 65288;
end
533:begin
x_i <= 65157;
end
534:begin
x_i <= 65160;
end
535:begin
x_i <= 65302;
end
536:begin
x_i <= 65330;
end
537:begin
x_i <= 65377;
end
538:begin
x_i <= 65485;
end
539:begin
x_i <= 55;
end
540:begin
x_i <= 131;
end
541:begin
x_i <= 86;
end
542:begin
x_i <= 103;
end
543:begin
x_i <= 87;
end
544:begin
x_i <= 105;
end
545:begin
x_i <= 57;
end
546:begin
x_i <= 40;
end
547:begin
x_i <= 6;
end
548:begin
x_i <= 65472;
end
549:begin
x_i <= 65469;
end
550:begin
x_i <= 65487;
end
551:begin
x_i <= 31;
end
552:begin
x_i <= 96;
end
553:begin
x_i <= 152;
end
554:begin
x_i <= 281;
end
555:begin
x_i <= 406;
end
556:begin
x_i <= 482;
end
557:begin
x_i <= 416;
end
558:begin
x_i <= 392;
end
559:begin
x_i <= 412;
end
560:begin
x_i <= 416;
end
561:begin
x_i <= 411;
end
562:begin
x_i <= 324;
end
563:begin
x_i <= 65307;
end
564:begin
x_i <= 64567;
end
565:begin
x_i <= 64488;
end
566:begin
x_i <= 64932;
end
567:begin
x_i <= 65478;
end
568:begin
x_i <= 61;
end
569:begin
x_i <= 136;
end
570:begin
x_i <= 597;
end
571:begin
x_i <= 672;
end
572:begin
x_i <= 354;
end
573:begin
x_i <= 210;
end
574:begin
x_i <= 83;
end
575:begin
x_i <= 65362;
end
576:begin
x_i <= 64911;
end
577:begin
x_i <= 64842;
end
578:begin
x_i <= 65330;
end
579:begin
x_i <= 12;
end
580:begin
x_i <= 19;
end
581:begin
x_i <= 143;
end
582:begin
x_i <= 367;
end
583:begin
x_i <= 282;
end
584:begin
x_i <= 13;
end
585:begin
x_i <= 65422;
end
586:begin
x_i <= 65409;
end
587:begin
x_i <= 65338;
end
588:begin
x_i <= 65204;
end
589:begin
x_i <= 65330;
end
590:begin
x_i <= 58;
end
591:begin
x_i <= 169;
end
592:begin
x_i <= 52;
end
593:begin
x_i <= 65479;
end
594:begin
x_i <= 65383;
end
595:begin
x_i <= 65190;
end
596:begin
x_i <= 65019;
end
597:begin
x_i <= 65048;
end
598:begin
x_i <= 65224;
end
599:begin
x_i <= 65348;
end
600:begin
x_i <= 65402;
end
601:begin
x_i <= 61;
end
602:begin
x_i <= 172;
end
603:begin
x_i <= 184;
end
604:begin
x_i <= 138;
end
605:begin
x_i <= 45;
end
606:begin
x_i <= 65472;
end
607:begin
x_i <= 65275;
end
608:begin
x_i <= 65195;
end
609:begin
x_i <= 65266;
end
610:begin
x_i <= 65287;
end
611:begin
x_i <= 65270;
end
612:begin
x_i <= 65348;
end
613:begin
x_i <= 65407;
end
614:begin
x_i <= 65474;
end
615:begin
x_i <= 18;
end
616:begin
x_i <= 91;
end
617:begin
x_i <= 135;
end
618:begin
x_i <= 245;
end
619:begin
x_i <= 202;
end
620:begin
x_i <= 163;
end
621:begin
x_i <= 104;
end
622:begin
x_i <= 65512;
end
623:begin
x_i <= 65448;
end
624:begin
x_i <= 65438;
end
625:begin
x_i <= 65476;
end
626:begin
x_i <= 65531;
end
627:begin
x_i <= 41;
end
628:begin
x_i <= 182;
end
629:begin
x_i <= 315;
end
630:begin
x_i <= 403;
end
631:begin
x_i <= 359;
end
632:begin
x_i <= 208;
end
633:begin
x_i <= 293;
end
634:begin
x_i <= 321;
end
635:begin
x_i <= 386;
end
636:begin
x_i <= 509;
end
637:begin
x_i <= 402;
end
638:begin
x_i <= 65478;
end
639:begin
x_i <= 64788;
end
640:begin
x_i <= 64712;
end
641:begin
x_i <= 65068;
end
642:begin
x_i <= 65384;
end
643:begin
x_i <= 65428;
end
644:begin
x_i <= 139;
end
645:begin
x_i <= 520;
end
646:begin
x_i <= 513;
end
647:begin
x_i <= 387;
end
648:begin
x_i <= 297;
end
649:begin
x_i <= 174;
end
650:begin
x_i <= 65366;
end
651:begin
x_i <= 65070;
end
652:begin
x_i <= 65088;
end
653:begin
x_i <= 65306;
end
654:begin
x_i <= 65437;
end
655:begin
x_i <= 65490;
end
656:begin
x_i <= 160;
end
657:begin
x_i <= 236;
end
658:begin
x_i <= 131;
end
659:begin
x_i <= 65535;
end
660:begin
x_i <= 65463;
end
661:begin
x_i <= 65427;
end
662:begin
x_i <= 65298;
end
663:begin
x_i <= 65219;
end
664:begin
x_i <= 65345;
end
665:begin
x_i <= 23;
end
666:begin
x_i <= 67;
end
667:begin
x_i <= 53;
end
668:begin
x_i <= 65514;
end
669:begin
x_i <= 65415;
end
670:begin
x_i <= 65348;
end
671:begin
x_i <= 65286;
end
672:begin
x_i <= 65253;
end
673:begin
x_i <= 65122;
end
674:begin
x_i <= 65034;
end
675:begin
x_i <= 65170;
end
676:begin
x_i <= 65316;
end
677:begin
x_i <= 65416;
end
678:begin
x_i <= 72;
end
679:begin
x_i <= 243;
end
680:begin
x_i <= 276;
end
681:begin
x_i <= 124;
end
682:begin
x_i <= 65502;
end
683:begin
x_i <= 65399;
end
684:begin
x_i <= 65214;
end
685:begin
x_i <= 65116;
end
686:begin
x_i <= 65099;
end
687:begin
x_i <= 65159;
end
688:begin
x_i <= 65306;
end
689:begin
x_i <= 65457;
end
690:begin
x_i <= 49;
end
691:begin
x_i <= 232;
end
692:begin
x_i <= 233;
end
693:begin
x_i <= 270;
end
694:begin
x_i <= 214;
end
695:begin
x_i <= 110;
end
696:begin
x_i <= 9;
end
697:begin
x_i <= 65444;
end
698:begin
x_i <= 65460;
end
699:begin
x_i <= 65478;
end
700:begin
x_i <= 65487;
end
701:begin
x_i <= 65527;
end
702:begin
x_i <= 70;
end
703:begin
x_i <= 247;
end
704:begin
x_i <= 299;
end
705:begin
x_i <= 450;
end
706:begin
x_i <= 562;
end
707:begin
x_i <= 666;
end
708:begin
x_i <= 738;
end
709:begin
x_i <= 745;
end
710:begin
x_i <= 725;
end
711:begin
x_i <= 25;
end
712:begin
x_i <= 64302;
end
713:begin
x_i <= 63845;
end
714:begin
x_i <= 64238;
end
715:begin
x_i <= 65104;
end
716:begin
x_i <= 0;
end
717:begin
x_i <= 125;
end
718:begin
x_i <= 849;
end
719:begin
x_i <= 1231;
end
720:begin
x_i <= 841;
end
721:begin
x_i <= 402;
end
722:begin
x_i <= 71;
end
723:begin
x_i <= 65160;
end
724:begin
x_i <= 64548;
end
725:begin
x_i <= 64337;
end
726:begin
x_i <= 64878;
end
727:begin
x_i <= 54;
end
728:begin
x_i <= 300;
end
729:begin
x_i <= 553;
end
730:begin
x_i <= 780;
end
731:begin
x_i <= 633;
end
732:begin
x_i <= 228;
end
733:begin
x_i <= 65281;
end
734:begin
x_i <= 65043;
end
735:begin
x_i <= 64930;
end
736:begin
x_i <= 64846;
end
737:begin
x_i <= 65052;
end
738:begin
x_i <= 35;
end
739:begin
x_i <= 395;
end
740:begin
x_i <= 466;
end
741:begin
x_i <= 346;
end
742:begin
x_i <= 175;
end
743:begin
x_i <= 65415;
end
744:begin
x_i <= 64986;
end
745:begin
x_i <= 64792;
end
746:begin
x_i <= 64845;
end
747:begin
x_i <= 65003;
end
748:begin
x_i <= 65193;
end
749:begin
x_i <= 65464;
end
750:begin
x_i <= 231;
end
751:begin
x_i <= 276;
end
752:begin
x_i <= 325;
end
753:begin
x_i <= 299;
end
754:begin
x_i <= 94;
end
755:begin
x_i <= 65418;
end
756:begin
x_i <= 65151;
end
757:begin
x_i <= 65135;
end
758:begin
x_i <= 65208;
end
759:begin
x_i <= 65138;
end
760:begin
x_i <= 65193;
end
761:begin
x_i <= 65287;
end
762:begin
x_i <= 65353;
end
763:begin
x_i <= 65528;
end
764:begin
x_i <= 81;
end
765:begin
x_i <= 139;
end
766:begin
x_i <= 299;
end
767:begin
x_i <= 337;
end
768:begin
x_i <= 288;
end
769:begin
x_i <= 178;
end
770:begin
x_i <= 16;
end
771:begin
x_i <= 65427;
end
772:begin
x_i <= 65347;
end
773:begin
x_i <= 65326;
end
774:begin
x_i <= 65362;
end
775:begin
x_i <= 65486;
end
776:begin
x_i <= 107;
end
777:begin
x_i <= 237;
end
778:begin
x_i <= 414;
end
779:begin
x_i <= 543;
end
780:begin
x_i <= 477;
end
781:begin
x_i <= 466;
end
782:begin
x_i <= 499;
end
783:begin
x_i <= 496;
end
784:begin
x_i <= 734;
end
785:begin
x_i <= 730;
end
786:begin
x_i <= 65495;
end
787:begin
x_i <= 64533;
end
788:begin
x_i <= 64140;
end
789:begin
x_i <= 64580;
end
790:begin
x_i <= 65225;
end
791:begin
x_i <= 65294;
end
792:begin
x_i <= 28;
end
793:begin
x_i <= 683;
end
794:begin
x_i <= 849;
end
795:begin
x_i <= 677;
end
796:begin
x_i <= 450;
end
797:begin
x_i <= 263;
end
798:begin
x_i <= 65406;
end
799:begin
x_i <= 64772;
end
800:begin
x_i <= 64608;
end
801:begin
x_i <= 65065;
end
802:begin
x_i <= 65443;
end
803:begin
x_i <= 78;
end
804:begin
x_i <= 379;
end
805:begin
x_i <= 560;
end
806:begin
x_i <= 454;
end
807:begin
x_i <= 88;
end
808:begin
x_i <= 65410;
end
809:begin
x_i <= 65290;
end
810:begin
x_i <= 65105;
end
811:begin
x_i <= 64913;
end
812:begin
x_i <= 65076;
end
813:begin
x_i <= 1;
end
814:begin
x_i <= 293;
end
815:begin
x_i <= 297;
end
816:begin
x_i <= 230;
end
817:begin
x_i <= 110;
end
818:begin
x_i <= 65402;
end
819:begin
x_i <= 65145;
end
820:begin
x_i <= 64937;
end
821:begin
x_i <= 64825;
end
822:begin
x_i <= 64758;
end
823:begin
x_i <= 64983;
end
824:begin
x_i <= 65368;
end
825:begin
x_i <= 206;
end
826:begin
x_i <= 390;
end
827:begin
x_i <= 430;
end
828:begin
x_i <= 348;
end
829:begin
x_i <= 190;
end
830:begin
x_i <= 65365;
end
831:begin
x_i <= 65161;
end
832:begin
x_i <= 65092;
end
833:begin
x_i <= 65041;
end
834:begin
x_i <= 65105;
end
835:begin
x_i <= 65215;
end
836:begin
x_i <= 65402;
end
837:begin
x_i <= 52;
end
838:begin
x_i <= 86;
end
839:begin
x_i <= 175;
end
840:begin
x_i <= 260;
end
841:begin
x_i <= 254;
end
842:begin
x_i <= 204;
end
843:begin
x_i <= 172;
end
844:begin
x_i <= 116;
end
845:begin
x_i <= 60;
end
846:begin
x_i <= 65520;
end
847:begin
x_i <= 65479;
end
848:begin
x_i <= 65476;
end
849:begin
x_i <= 12;
end
850:begin
x_i <= 79;
end
851:begin
x_i <= 225;
end
852:begin
x_i <= 419;
end
853:begin
x_i <= 556;
end
854:begin
x_i <= 693;
end
855:begin
x_i <= 707;
end
856:begin
x_i <= 800;
end
857:begin
x_i <= 1059;
end
858:begin
x_i <= 828;
end
859:begin
x_i <= 65011;
end
860:begin
x_i <= 63667;
end
861:begin
x_i <= 63589;
end
862:begin
x_i <= 64502;
end
863:begin
x_i <= 65332;
end
864:begin
x_i <= 65465;
end
865:begin
x_i <= 460;
end
866:begin
x_i <= 1318;
end
867:begin
x_i <= 1271;
end
868:begin
x_i <= 783;
end
869:begin
x_i <= 433;
end
870:begin
x_i <= 1;
end
871:begin
x_i <= 64781;
end
872:begin
x_i <= 64088;
end
873:begin
x_i <= 64285;
end
874:begin
x_i <= 65186;
end
875:begin
x_i <= 235;
end
876:begin
x_i <= 513;
end
877:begin
x_i <= 908;
end
878:begin
x_i <= 949;
end
879:begin
x_i <= 564;
end
880:begin
x_i <= 47;
end
881:begin
x_i <= 65183;
end
882:begin
x_i <= 64908;
end
883:begin
x_i <= 64641;
end
884:begin
x_i <= 64659;
end
885:begin
x_i <= 65237;
end
886:begin
x_i <= 291;
end
887:begin
x_i <= 557;
end
888:begin
x_i <= 552;
end
889:begin
x_i <= 398;
end
890:begin
x_i <= 85;
end
891:begin
x_i <= 65175;
end
892:begin
x_i <= 64857;
end
893:begin
x_i <= 64728;
end
894:begin
x_i <= 64656;
end
895:begin
x_i <= 64675;
end
896:begin
x_i <= 65043;
end
897:begin
x_i <= 25;
end
898:begin
x_i <= 376;
end
899:begin
x_i <= 600;
end
900:begin
x_i <= 696;
end
901:begin
x_i <= 566;
end
902:begin
x_i <= 92;
end
903:begin
x_i <= 65193;
end
904:begin
x_i <= 65014;
end
905:begin
x_i <= 64985;
end
906:begin
x_i <= 64933;
end
907:begin
x_i <= 65028;
end
908:begin
x_i <= 65270;
end
909:begin
x_i <= 65496;
end
910:begin
x_i <= 170;
end
911:begin
x_i <= 317;
end
912:begin
x_i <= 371;
end
913:begin
x_i <= 343;
end
914:begin
x_i <= 275;
end
915:begin
x_i <= 248;
end
916:begin
x_i <= 205;
end
917:begin
x_i <= 44;
end
918:begin
x_i <= 65437;
end
919:begin
x_i <= 65424;
end
920:begin
x_i <= 65433;
end
921:begin
x_i <= 65527;
end
922:begin
x_i <= 100;
end
923:begin
x_i <= 262;
end
924:begin
x_i <= 436;
end
925:begin
x_i <= 545;
end
926:begin
x_i <= 779;
end
927:begin
x_i <= 874;
end
928:begin
x_i <= 905;
end
929:begin
x_i <= 988;
end
930:begin
x_i <= 813;
end
931:begin
x_i <= 65006;
end
932:begin
x_i <= 63589;
end
933:begin
x_i <= 63477;
end
934:begin
x_i <= 64411;
end
935:begin
x_i <= 65387;
end
936:begin
x_i <= 65513;
end
937:begin
x_i <= 528;
end
938:begin
x_i <= 1400;
end
939:begin
x_i <= 1289;
end
940:begin
x_i <= 730;
end
941:begin
x_i <= 430;
end
942:begin
x_i <= 64;
end
943:begin
x_i <= 64778;
end
944:begin
x_i <= 63996;
end
945:begin
x_i <= 64203;
end
946:begin
x_i <= 65160;
end
947:begin
x_i <= 240;
end
948:begin
x_i <= 538;
end
949:begin
x_i <= 974;
end
950:begin
x_i <= 1041;
end
951:begin
x_i <= 614;
end
952:begin
x_i <= 82;
end
953:begin
x_i <= 65224;
end
954:begin
x_i <= 64932;
end
955:begin
x_i <= 64566;
end
956:begin
x_i <= 64505;
end
957:begin
x_i <= 65107;
end
958:begin
x_i <= 369;
end
959:begin
x_i <= 672;
end
960:begin
x_i <= 604;
end
961:begin
x_i <= 460;
end
962:begin
x_i <= 104;
end
963:begin
x_i <= 65146;
end
964:begin
x_i <= 64789;
end
965:begin
x_i <= 64733;
end
966:begin
x_i <= 64723;
end
967:begin
x_i <= 64717;
end
968:begin
x_i <= 65058;
end
969:begin
x_i <= 77;
end
970:begin
x_i <= 444;
end
971:begin
x_i <= 569;
end
972:begin
x_i <= 605;
end
973:begin
x_i <= 442;
end
974:begin
x_i <= 65525;
end
975:begin
x_i <= 65075;
end
976:begin
x_i <= 64937;
end
977:begin
x_i <= 65002;
end
978:begin
x_i <= 64986;
end
979:begin
x_i <= 65065;
end
980:begin
x_i <= 65291;
end
981:begin
x_i <= 14;
end
982:begin
x_i <= 196;
end
983:begin
x_i <= 318;
end
984:begin
x_i <= 394;
end
985:begin
x_i <= 363;
end
986:begin
x_i <= 301;
end
987:begin
x_i <= 269;
end
988:begin
x_i <= 209;
end
989:begin
x_i <= 64;
end
990:begin
x_i <= 65463;
end
991:begin
x_i <= 65389;
end
992:begin
x_i <= 65409;
end
993:begin
x_i <= 3;
end
994:begin
x_i <= 135;
end
995:begin
x_i <= 399;
end
996:begin
x_i <= 547;
end
997:begin
x_i <= 707;
end
998:begin
x_i <= 920;
end
999:begin
x_i <= 1018;
end
1000:begin
x_i <= 1065;
end
1001:begin
x_i <= 1023;
end
1002:begin
x_i <= 113;
end
1003:begin
x_i <= 64074;
end
1004:begin
x_i <= 63398;
end
1005:begin
x_i <= 63841;
end
1006:begin
x_i <= 64868;
end
1007:begin
x_i <= 65459;
end
1008:begin
x_i <= 229;
end
1009:begin
x_i <= 1173;
end
1010:begin
x_i <= 1565;
end
1011:begin
x_i <= 984;
end
1012:begin
x_i <= 591;
end
1013:begin
x_i <= 260;
end
1014:begin
x_i <= 65119;
end
1015:begin
x_i <= 64277;
end
1016:begin
x_i <= 64041;
end
1017:begin
x_i <= 64770;
end
1018:begin
x_i <= 3;
end
1019:begin
x_i <= 331;
end
1020:begin
x_i <= 848;
end
1021:begin
x_i <= 1182;
end
1022:begin
x_i <= 868;
end
1023:begin
x_i <= 275;
end
1024:begin
x_i <= 65359;
end
1025:begin
x_i <= 65098;
end
1026:begin
x_i <= 64773;
end
1027:begin
x_i <= 64467;
end
1028:begin
x_i <= 64804;
end
1029:begin
x_i <= 27;
end
1030:begin
x_i <= 536;
end
1031:begin
x_i <= 602;
end
1032:begin
x_i <= 587;
end
1033:begin
x_i <= 446;
end
1034:begin
x_i <= 60;
end
1035:begin
x_i <= 65042;
end
1036:begin
x_i <= 64637;
end
1037:begin
x_i <= 64575;
end
1038:begin
x_i <= 64616;
end
1039:begin
x_i <= 64885;
end
1040:begin
x_i <= 65350;
end
1041:begin
x_i <= 363;
end
1042:begin
x_i <= 684;
end
1043:begin
x_i <= 740;
end
1044:begin
x_i <= 474;
end
1045:begin
x_i <= 72;
end
1046:begin
x_i <= 65119;
end
1047:begin
x_i <= 64828;
end
1048:begin
x_i <= 64846;
end
1049:begin
x_i <= 64909;
end
1050:begin
x_i <= 65098;
end
1051:begin
x_i <= 65265;
end
1052:begin
x_i <= 65450;
end
1053:begin
x_i <= 114;
end
1054:begin
x_i <= 221;
end
1055:begin
x_i <= 254;
end
1056:begin
x_i <= 242;
end
1057:begin
x_i <= 188;
end
1058:begin
x_i <= 242;
end
1059:begin
x_i <= 239;
end
1060:begin
x_i <= 206;
end
1061:begin
x_i <= 166;
end
1062:begin
x_i <= 73;
end
1063:begin
x_i <= 65491;
end
1064:begin
x_i <= 65444;
end
1065:begin
x_i <= 65484;
end
1066:begin
x_i <= 110;
end
1067:begin
x_i <= 314;
end
1068:begin
x_i <= 462;
end
1069:begin
x_i <= 733;
end
1070:begin
x_i <= 1017;
end
1071:begin
x_i <= 1124;
end
1072:begin
x_i <= 976;
end
1073:begin
x_i <= 753;
end
1074:begin
x_i <= 304;
end
1075:begin
x_i <= 64528;
end
1076:begin
x_i <= 63518;
end
1077:begin
x_i <= 63661;
end
1078:begin
x_i <= 64570;
end
1079:begin
x_i <= 65501;
end
1080:begin
x_i <= 272;
end
1081:begin
x_i <= 917;
end
1082:begin
x_i <= 1625;
end
1083:begin
x_i <= 1235;
end
1084:begin
x_i <= 591;
end
1085:begin
x_i <= 166;
end
1086:begin
x_i <= 65181;
end
1087:begin
x_i <= 64513;
end
1088:begin
x_i <= 64105;
end
1089:begin
x_i <= 64516;
end
1090:begin
x_i <= 65433;
end
1091:begin
x_i <= 429;
end
1092:begin
x_i <= 749;
end
1093:begin
x_i <= 1096;
end
1094:begin
x_i <= 916;
end
1095:begin
x_i <= 368;
end
1096:begin
x_i <= 65384;
end
1097:begin
x_i <= 65012;
end
1098:begin
x_i <= 64806;
end
1099:begin
x_i <= 64634;
end
1100:begin
x_i <= 64841;
end
1101:begin
x_i <= 65440;
end
1102:begin
x_i <= 462;
end
1103:begin
x_i <= 625;
end
1104:begin
x_i <= 493;
end
1105:begin
x_i <= 205;
end
1106:begin
x_i <= 65392;
end
1107:begin
x_i <= 65016;
end
1108:begin
x_i <= 64798;
end
1109:begin
x_i <= 64773;
end
1110:begin
x_i <= 64878;
end
1111:begin
x_i <= 65006;
end
1112:begin
x_i <= 65286;
end
1113:begin
x_i <= 88;
end
1114:begin
x_i <= 432;
end
1115:begin
x_i <= 518;
end
1116:begin
x_i <= 470;
end
1117:begin
x_i <= 244;
end
1118:begin
x_i <= 65409;
end
1119:begin
x_i <= 65090;
end
1120:begin
x_i <= 64953;
end
1121:begin
x_i <= 64913;
end
1122:begin
x_i <= 65039;
end
1123:begin
x_i <= 65155;
end
1124:begin
x_i <= 65269;
end
1125:begin
x_i <= 65515;
end
1126:begin
x_i <= 179;
end
1127:begin
x_i <= 321;
end
1128:begin
x_i <= 411;
end
1129:begin
x_i <= 414;
end
1130:begin
x_i <= 401;
end
1131:begin
x_i <= 366;
end
1132:begin
x_i <= 230;
end
1133:begin
x_i <= 87;
end
1134:begin
x_i <= 65479;
end
1135:begin
x_i <= 65439;
end
1136:begin
x_i <= 65508;
end
1137:begin
x_i <= 74;
end
1138:begin
x_i <= 330;
end
1139:begin
x_i <= 587;
end
1140:begin
x_i <= 851;
end
1141:begin
x_i <= 1084;
end
1142:begin
x_i <= 1223;
end
1143:begin
x_i <= 1122;
end
1144:begin
x_i <= 765;
end
1145:begin
x_i <= 64847;
end
1146:begin
x_i <= 63493;
end
1147:begin
x_i <= 63495;
end
1148:begin
x_i <= 64200;
end
1149:begin
x_i <= 65103;
end
1150:begin
x_i <= 40;
end
1151:begin
x_i <= 781;
end
1152:begin
x_i <= 1720;
end
1153:begin
x_i <= 1507;
end
1154:begin
x_i <= 801;
end
1155:begin
x_i <= 524;
end
1156:begin
x_i <= 65469;
end
1157:begin
x_i <= 64496;
end
1158:begin
x_i <= 63891;
end
1159:begin
x_i <= 64250;
end
1160:begin
x_i <= 65166;
end
1161:begin
x_i <= 268;
end
1162:begin
x_i <= 620;
end
1163:begin
x_i <= 1172;
end
1164:begin
x_i <= 1153;
end
1165:begin
x_i <= 629;
end
1166:begin
x_i <= 49;
end
1167:begin
x_i <= 65171;
end
1168:begin
x_i <= 64833;
end
1169:begin
x_i <= 64535;
end
1170:begin
x_i <= 64592;
end
1171:begin
x_i <= 65162;
end
1172:begin
x_i <= 323;
end
1173:begin
x_i <= 650;
end
1174:begin
x_i <= 703;
end
1175:begin
x_i <= 438;
end
1176:begin
x_i <= 18;
end
1177:begin
x_i <= 65104;
end
1178:begin
x_i <= 64803;
end
1179:begin
x_i <= 64692;
end
1180:begin
x_i <= 64550;
end
1181:begin
x_i <= 64611;
end
1182:begin
x_i <= 65110;
end
1183:begin
x_i <= 164;
end
1184:begin
x_i <= 489;
end
1185:begin
x_i <= 659;
end
1186:begin
x_i <= 710;
end
1187:begin
x_i <= 534;
end
1188:begin
x_i <= 65513;
end
1189:begin
x_i <= 65053;
end
1190:begin
x_i <= 64940;
end
1191:begin
x_i <= 64859;
end
1192:begin
x_i <= 64766;
end
1193:begin
x_i <= 64921;
end
1194:begin
x_i <= 65244;
end
1195:begin
x_i <= 65517;
end
1196:begin
x_i <= 169;
end
1197:begin
x_i <= 327;
end
1198:begin
x_i <= 468;
end
1199:begin
x_i <= 476;
end
1200:begin
x_i <= 402;
end
1201:begin
x_i <= 417;
end
1202:begin
x_i <= 322;
end
1203:begin
x_i <= 169;
end
1204:begin
x_i <= 35;
end
1205:begin
x_i <= 65521;
end
1206:begin
x_i <= 67;
end
1207:begin
x_i <= 130;
end
1208:begin
x_i <= 302;
end
1209:begin
x_i <= 566;
end
1210:begin
x_i <= 840;
end
1211:begin
x_i <= 1020;
end
1212:begin
x_i <= 1093;
end
1213:begin
x_i <= 1132;
end
1214:begin
x_i <= 660;
end
1215:begin
x_i <= 64598;
end
1216:begin
x_i <= 63463;
end
1217:begin
x_i <= 63719;
end
1218:begin
x_i <= 64509;
end
1219:begin
x_i <= 65208;
end
1220:begin
x_i <= 65509;
end
1221:begin
x_i <= 874;
end
1222:begin
x_i <= 1715;
end
1223:begin
x_i <= 1226;
end
1224:begin
x_i <= 656;
end
1225:begin
x_i <= 486;
end
1226:begin
x_i <= 65384;
end
1227:begin
x_i <= 64345;
end
1228:begin
x_i <= 63826;
end
1229:begin
x_i <= 64408;
end
1230:begin
x_i <= 65396;
end
1231:begin
x_i <= 380;
end
1232:begin
x_i <= 715;
end
1233:begin
x_i <= 1272;
end
1234:begin
x_i <= 1135;
end
1235:begin
x_i <= 482;
end
1236:begin
x_i <= 65426;
end
1237:begin
x_i <= 65021;
end
1238:begin
x_i <= 64650;
end
1239:begin
x_i <= 64416;
end
1240:begin
x_i <= 64590;
end
1241:begin
x_i <= 65331;
end
1242:begin
x_i <= 533;
end
1243:begin
x_i <= 775;
end
1244:begin
x_i <= 734;
end
1245:begin
x_i <= 440;
end
1246:begin
x_i <= 65393;
end
1247:begin
x_i <= 64862;
end
1248:begin
x_i <= 64689;
end
1249:begin
x_i <= 64602;
end
1250:begin
x_i <= 64517;
end
1251:begin
x_i <= 64626;
end
1252:begin
x_i <= 65215;
end
1253:begin
x_i <= 365;
end
1254:begin
x_i <= 658;
end
1255:begin
x_i <= 702;
end
1256:begin
x_i <= 718;
end
1257:begin
x_i <= 437;
end
1258:begin
x_i <= 65383;
end
1259:begin
x_i <= 65009;
end
1260:begin
x_i <= 64889;
end
1261:begin
x_i <= 64842;
end
1262:begin
x_i <= 64841;
end
1263:begin
x_i <= 65036;
end
1264:begin
x_i <= 65350;
end
1265:begin
x_i <= 94;
end
1266:begin
x_i <= 239;
end
1267:begin
x_i <= 300;
end
1268:begin
x_i <= 364;
end
1269:begin
x_i <= 355;
end
1270:begin
x_i <= 346;
end
1271:begin
x_i <= 357;
end
1272:begin
x_i <= 290;
end
1273:begin
x_i <= 215;
end
1274:begin
x_i <= 103;
end
1275:begin
x_i <= 152;
end
1276:begin
x_i <= 239;
end
1277:begin
x_i <= 324;
end
1278:begin
x_i <= 491;
end
1279:begin
x_i <= 692;
end
1280:begin
x_i <= 862;
end
1281:begin
x_i <= 980;
end
1282:begin
x_i <= 988;
end
1283:begin
x_i <= 880;
end
1284:begin
x_i <= 65231;
end
1285:begin
x_i <= 63697;
end
1286:begin
x_i <= 63578;
end
1287:begin
x_i <= 64236;
end
1288:begin
x_i <= 64992;
end
1289:begin
x_i <= 65428;
end
1290:begin
x_i <= 538;
end
1291:begin
x_i <= 1493;
end
1292:begin
x_i <= 1348;
end
1293:begin
x_i <= 697;
end
1294:begin
x_i <= 545;
end
1295:begin
x_i <= 106;
end
1296:begin
x_i <= 64672;
end
1297:begin
x_i <= 63975;
end
1298:begin
x_i <= 64239;
end
1299:begin
x_i <= 65072;
end
1300:begin
x_i <= 158;
end
1301:begin
x_i <= 640;
end
1302:begin
x_i <= 1209;
end
1303:begin
x_i <= 1274;
end
1304:begin
x_i <= 632;
end
1305:begin
x_i <= 75;
end
1306:begin
x_i <= 65187;
end
1307:begin
x_i <= 64713;
end
1308:begin
x_i <= 64310;
end
1309:begin
x_i <= 64424;
end
1310:begin
x_i <= 65117;
end
1311:begin
x_i <= 317;
end
1312:begin
x_i <= 748;
end
1313:begin
x_i <= 848;
end
1314:begin
x_i <= 684;
end
1315:begin
x_i <= 193;
end
1316:begin
x_i <= 65068;
end
1317:begin
x_i <= 64829;
end
1318:begin
x_i <= 64775;
end
1319:begin
x_i <= 64528;
end
1320:begin
x_i <= 64418;
end
1321:begin
x_i <= 64765;
end
1322:begin
x_i <= 47;
end
1323:begin
x_i <= 517;
end
1324:begin
x_i <= 623;
end
1325:begin
x_i <= 823;
end
1326:begin
x_i <= 687;
end
1327:begin
x_i <= 148;
end
1328:begin
x_i <= 65196;
end
1329:begin
x_i <= 64949;
end
1330:begin
x_i <= 64863;
end
1331:begin
x_i <= 64683;
end
1332:begin
x_i <= 64787;
end
1333:begin
x_i <= 65175;
end
1334:begin
x_i <= 3;
end
1335:begin
x_i <= 206;
end
1336:begin
x_i <= 388;
end
1337:begin
x_i <= 500;
end
1338:begin
x_i <= 501;
end
1339:begin
x_i <= 399;
end
1340:begin
x_i <= 351;
end
1341:begin
x_i <= 238;
end
1342:begin
x_i <= 38;
end
1343:begin
x_i <= 65467;
end
1344:begin
x_i <= 16;
end
1345:begin
x_i <= 166;
end
1346:begin
x_i <= 369;
end
1347:begin
x_i <= 550;
end
1348:begin
x_i <= 813;
end
1349:begin
x_i <= 1045;
end
1350:begin
x_i <= 1005;
end
1351:begin
x_i <= 839;
end
1352:begin
x_i <= 830;
end
1353:begin
x_i <= 90;
end
1354:begin
x_i <= 64149;
end
1355:begin
x_i <= 63627;
end
1356:begin
x_i <= 64079;
end
1357:begin
x_i <= 64883;
end
1358:begin
x_i <= 65428;
end
1359:begin
x_i <= 246;
end
1360:begin
x_i <= 1308;
end
1361:begin
x_i <= 1468;
end
1362:begin
x_i <= 684;
end
1363:begin
x_i <= 385;
end
1364:begin
x_i <= 135;
end
1365:begin
x_i <= 64905;
end
1366:begin
x_i <= 64188;
end
1367:begin
x_i <= 64262;
end
1368:begin
x_i <= 65043;
end
1369:begin
x_i <= 158;
end
1370:begin
x_i <= 509;
end
1371:begin
x_i <= 1101;
end
1372:begin
x_i <= 1330;
end
1373:begin
x_i <= 734;
end
1374:begin
x_i <= 109;
end
1375:begin
x_i <= 65211;
end
1376:begin
x_i <= 64839;
end
1377:begin
x_i <= 64453;
end
1378:begin
x_i <= 64374;
end
1379:begin
x_i <= 64843;
end
1380:begin
x_i <= 44;
end
1381:begin
x_i <= 510;
end
1382:begin
x_i <= 714;
end
1383:begin
x_i <= 704;
end
1384:begin
x_i <= 397;
end
1385:begin
x_i <= 65342;
end
1386:begin
x_i <= 64764;
end
1387:begin
x_i <= 64673;
end
1388:begin
x_i <= 64619;
end
1389:begin
x_i <= 64606;
end
1390:begin
x_i <= 64967;
end
1391:begin
x_i <= 65531;
end
1392:begin
x_i <= 535;
end
1393:begin
x_i <= 658;
end
1394:begin
x_i <= 602;
end
1395:begin
x_i <= 520;
end
1396:begin
x_i <= 50;
end
1397:begin
x_i <= 65081;
end
1398:begin
x_i <= 64938;
end
1399:begin
x_i <= 64894;
end
1400:begin
x_i <= 64893;
end
1401:begin
x_i <= 65055;
end
1402:begin
x_i <= 65363;
end
1403:begin
x_i <= 66;
end
1404:begin
x_i <= 173;
end
1405:begin
x_i <= 244;
end
1406:begin
x_i <= 318;
end
1407:begin
x_i <= 250;
end
1408:begin
x_i <= 143;
end
1409:begin
x_i <= 210;
end
1410:begin
x_i <= 302;
end
1411:begin
x_i <= 237;
end
1412:begin
x_i <= 143;
end
1413:begin
x_i <= 153;
end
1414:begin
x_i <= 311;
end
1415:begin
x_i <= 384;
end
1416:begin
x_i <= 446;
end
1417:begin
x_i <= 592;
end
1418:begin
x_i <= 788;
end
1419:begin
x_i <= 908;
end
1420:begin
x_i <= 935;
end
1421:begin
x_i <= 1021;
end
1422:begin
x_i <= 394;
end
1423:begin
x_i <= 64430;
end
1424:begin
x_i <= 63724;
end
1425:begin
x_i <= 64188;
end
1426:begin
x_i <= 64836;
end
1427:begin
x_i <= 65218;
end
1428:begin
x_i <= 51;
end
1429:begin
x_i <= 1024;
end
1430:begin
x_i <= 1253;
end
1431:begin
x_i <= 548;
end
1432:begin
x_i <= 396;
end
1433:begin
x_i <= 333;
end
1434:begin
x_i <= 65074;
end
1435:begin
x_i <= 64244;
end
1436:begin
x_i <= 64359;
end
1437:begin
x_i <= 65113;
end
1438:begin
x_i <= 148;
end
1439:begin
x_i <= 489;
end
1440:begin
x_i <= 1038;
end
1441:begin
x_i <= 1295;
end
1442:begin
x_i <= 702;
end
1443:begin
x_i <= 46;
end
1444:begin
x_i <= 65296;
end
1445:begin
x_i <= 64895;
end
1446:begin
x_i <= 64449;
end
1447:begin
x_i <= 64351;
end
1448:begin
x_i <= 64852;
end
1449:begin
x_i <= 47;
end
1450:begin
x_i <= 431;
end
1451:begin
x_i <= 674;
end
1452:begin
x_i <= 620;
end
1453:begin
x_i <= 243;
end
1454:begin
x_i <= 65216;
end
1455:begin
x_i <= 64808;
end
1456:begin
x_i <= 64629;
end
1457:begin
x_i <= 64536;
end
1458:begin
x_i <= 64535;
end
1459:begin
x_i <= 65007;
end
1460:begin
x_i <= 181;
end
1461:begin
x_i <= 618;
end
1462:begin
x_i <= 775;
end
1463:begin
x_i <= 791;
end
1464:begin
x_i <= 563;
end
1465:begin
x_i <= 31;
end
1466:begin
x_i <= 65035;
end
1467:begin
x_i <= 64872;
end
1468:begin
x_i <= 64743;
end
1469:begin
x_i <= 64782;
end
1470:begin
x_i <= 65077;
end
1471:begin
x_i <= 65482;
end
1472:begin
x_i <= 260;
end
1473:begin
x_i <= 361;
end
1474:begin
x_i <= 437;
end
1475:begin
x_i <= 421;
end
1476:begin
x_i <= 176;
end
1477:begin
x_i <= 18;
end
1478:begin
x_i <= 63;
end
1479:begin
x_i <= 118;
end
1480:begin
x_i <= 91;
end
1481:begin
x_i <= 183;
end
1482:begin
x_i <= 415;
end
1483:begin
x_i <= 567;
end
1484:begin
x_i <= 598;
end
1485:begin
x_i <= 585;
end
1486:begin
x_i <= 650;
end
1487:begin
x_i <= 774;
end
1488:begin
x_i <= 725;
end
1489:begin
x_i <= 832;
end
1490:begin
x_i <= 887;
end
1491:begin
x_i <= 65403;
end
1492:begin
x_i <= 64182;
end
1493:begin
x_i <= 64046;
end
1494:begin
x_i <= 64591;
end
1495:begin
x_i <= 65150;
end
1496:begin
x_i <= 65316;
end
1497:begin
x_i <= 379;
end
1498:begin
x_i <= 1142;
end
1499:begin
x_i <= 763;
end
1500:begin
x_i <= 280;
end
1501:begin
x_i <= 410;
end
1502:begin
x_i <= 24;
end
1503:begin
x_i <= 64661;
end
1504:begin
x_i <= 64219;
end
1505:begin
x_i <= 64702;
end
1506:begin
x_i <= 65352;
end
1507:begin
x_i <= 152;
end
1508:begin
x_i <= 707;
end
1509:begin
x_i <= 1331;
end
1510:begin
x_i <= 1090;
end
1511:begin
x_i <= 403;
end
1512:begin
x_i <= 32;
end
1513:begin
x_i <= 65257;
end
1514:begin
x_i <= 64730;
end
1515:begin
x_i <= 64334;
end
1516:begin
x_i <= 64502;
end
1517:begin
x_i <= 65094;
end
1518:begin
x_i <= 41;
end
1519:begin
x_i <= 401;
end
1520:begin
x_i <= 578;
end
1521:begin
x_i <= 423;
end
1522:begin
x_i <= 65500;
end
1523:begin
x_i <= 65040;
end
1524:begin
x_i <= 64798;
end
1525:begin
x_i <= 64658;
end
1526:begin
x_i <= 64478;
end
1527:begin
x_i <= 64666;
end
1528:begin
x_i <= 65173;
end
1529:begin
x_i <= 289;
end
1530:begin
x_i <= 650;
end
1531:begin
x_i <= 751;
end
1532:begin
x_i <= 850;
end
1533:begin
x_i <= 499;
end
1534:begin
x_i <= 65427;
end
1535:begin
x_i <= 65097;
end
1536:begin
x_i <= 64921;
end
1537:begin
x_i <= 64857;
end
1538:begin
x_i <= 64870;
end
1539:begin
x_i <= 65094;
end
1540:begin
x_i <= 65490;
end
1541:begin
x_i <= 169;
end
1542:begin
x_i <= 351;
end
1543:begin
x_i <= 490;
end
1544:begin
x_i <= 387;
end
1545:begin
x_i <= 190;
end
1546:begin
x_i <= 112;
end
1547:begin
x_i <= 170;
end
1548:begin
x_i <= 185;
end
1549:begin
x_i <= 132;
end
1550:begin
x_i <= 218;
end
1551:begin
x_i <= 412;
end
1552:begin
x_i <= 570;
end
1553:begin
x_i <= 668;
end
1554:begin
x_i <= 732;
end
1555:begin
x_i <= 770;
end
1556:begin
x_i <= 812;
end
1557:begin
x_i <= 900;
end
1558:begin
x_i <= 956;
end
1559:begin
x_i <= 65404;
end
1560:begin
x_i <= 64229;
end
1561:begin
x_i <= 64070;
end
1562:begin
x_i <= 64511;
end
1563:begin
x_i <= 65097;
end
1564:begin
x_i <= 65336;
end
1565:begin
x_i <= 438;
end
1566:begin
x_i <= 1083;
end
1567:begin
x_i <= 560;
end
1568:begin
x_i <= 181;
end
1569:begin
x_i <= 444;
end
1570:begin
x_i <= 94;
end
1571:begin
x_i <= 64695;
end
1572:begin
x_i <= 64275;
end
1573:begin
x_i <= 64781;
end
1574:begin
x_i <= 65350;
end
1575:begin
x_i <= 22;
end
1576:begin
x_i <= 554;
end
1577:begin
x_i <= 1286;
end
1578:begin
x_i <= 1046;
end
1579:begin
x_i <= 339;
end
1580:begin
x_i <= 121;
end
1581:begin
x_i <= 65439;
end
1582:begin
x_i <= 64923;
end
1583:begin
x_i <= 64454;
end
1584:begin
x_i <= 64567;
end
1585:begin
x_i <= 65119;
end
1586:begin
x_i <= 65463;
end
1587:begin
x_i <= 298;
end
1588:begin
x_i <= 565;
end
1589:begin
x_i <= 369;
end
1590:begin
x_i <= 65434;
end
1591:begin
x_i <= 64987;
end
1592:begin
x_i <= 64754;
end
1593:begin
x_i <= 64595;
end
1594:begin
x_i <= 64437;
end
1595:begin
x_i <= 64636;
end
1596:begin
x_i <= 65141;
end
1597:begin
x_i <= 189;
end
1598:begin
x_i <= 525;
end
1599:begin
x_i <= 733;
end
1600:begin
x_i <= 814;
end
1601:begin
x_i <= 541;
end
1602:begin
x_i <= 65482;
end
1603:begin
x_i <= 65095;
end
1604:begin
x_i <= 64992;
end
1605:begin
x_i <= 64917;
end
1606:begin
x_i <= 64923;
end
1607:begin
x_i <= 65223;
end
1608:begin
x_i <= 10;
end
1609:begin
x_i <= 151;
end
1610:begin
x_i <= 281;
end
1611:begin
x_i <= 387;
end
1612:begin
x_i <= 294;
end
1613:begin
x_i <= 34;
end
1614:begin
x_i <= 12;
end
1615:begin
x_i <= 131;
end
1616:begin
x_i <= 170;
end
1617:begin
x_i <= 224;
end
1618:begin
x_i <= 407;
end
1619:begin
x_i <= 611;
end
1620:begin
x_i <= 661;
end
1621:begin
x_i <= 627;
end
1622:begin
x_i <= 643;
end
1623:begin
x_i <= 692;
end
1624:begin
x_i <= 628;
end
1625:begin
x_i <= 873;
end
1626:begin
x_i <= 927;
end
1627:begin
x_i <= 65457;
end
1628:begin
x_i <= 64426;
end
1629:begin
x_i <= 64366;
end
1630:begin
x_i <= 64806;
end
1631:begin
x_i <= 65108;
end
1632:begin
x_i <= 65123;
end
1633:begin
x_i <= 301;
end
1634:begin
x_i <= 826;
end
1635:begin
x_i <= 286;
end
1636:begin
x_i <= 141;
end
1637:begin
x_i <= 395;
end
1638:begin
x_i <= 107;
end
1639:begin
x_i <= 64789;
end
1640:begin
x_i <= 64363;
end
1641:begin
x_i <= 65015;
end
1642:begin
x_i <= 65405;
end
1643:begin
x_i <= 65481;
end
1644:begin
x_i <= 529;
end
1645:begin
x_i <= 1118;
end
1646:begin
x_i <= 851;
end
1647:begin
x_i <= 354;
end
1648:begin
x_i <= 249;
end
1649:begin
x_i <= 100;
end
1650:begin
x_i <= 65028;
end
1651:begin
x_i <= 64531;
end
1652:begin
x_i <= 64724;
end
1653:begin
x_i <= 65083;
end
1654:begin
x_i <= 65326;
end
1655:begin
x_i <= 85;
end
1656:begin
x_i <= 344;
end
1657:begin
x_i <= 184;
end
1658:begin
x_i <= 65386;
end
1659:begin
x_i <= 65065;
end
1660:begin
x_i <= 64908;
end
1661:begin
x_i <= 64682;
end
1662:begin
x_i <= 64454;
end
1663:begin
x_i <= 64758;
end
1664:begin
x_i <= 65150;
end
1665:begin
x_i <= 77;
end
1666:begin
x_i <= 460;
end
1667:begin
x_i <= 539;
end
1668:begin
x_i <= 698;
end
1669:begin
x_i <= 454;
end
1670:begin
x_i <= 33;
end
1671:begin
x_i <= 65296;
end
1672:begin
x_i <= 65143;
end
1673:begin
x_i <= 65075;
end
1674:begin
x_i <= 65107;
end
1675:begin
x_i <= 65300;
end
1676:begin
x_i <= 74;
end
1677:begin
x_i <= 201;
end
1678:begin
x_i <= 268;
end
1679:begin
x_i <= 322;
end
1680:begin
x_i <= 231;
end
1681:begin
x_i <= 5;
end
1682:begin
x_i <= 65513;
end
1683:begin
x_i <= 84;
end
1684:begin
x_i <= 28;
end
1685:begin
x_i <= 124;
end
1686:begin
x_i <= 418;
end
1687:begin
x_i <= 636;
end
1688:begin
x_i <= 682;
end
1689:begin
x_i <= 649;
end
1690:begin
x_i <= 684;
end
1691:begin
x_i <= 660;
end
1692:begin
x_i <= 540;
end
1693:begin
x_i <= 722;
end
1694:begin
x_i <= 862;
end
1695:begin
x_i <= 68;
end
1696:begin
x_i <= 64758;
end
1697:begin
x_i <= 64697;
end
1698:begin
x_i <= 64991;
end
1699:begin
x_i <= 65290;
end
1700:begin
x_i <= 65368;
end
1701:begin
x_i <= 177;
end
1702:begin
x_i <= 362;
end
1703:begin
x_i <= 65505;
end
1704:begin
x_i <= 65450;
end
1705:begin
x_i <= 181;
end
1706:begin
x_i <= 30;
end
1707:begin
x_i <= 65054;
end
1708:begin
x_i <= 64810;
end
1709:begin
x_i <= 65060;
end
1710:begin
x_i <= 65290;
end
1711:begin
x_i <= 65506;
end
1712:begin
x_i <= 382;
end
1713:begin
x_i <= 689;
end
1714:begin
x_i <= 583;
end
1715:begin
x_i <= 348;
end
1716:begin
x_i <= 353;
end
1717:begin
x_i <= 248;
end
1718:begin
x_i <= 65441;
end
1719:begin
x_i <= 65110;
end
1720:begin
x_i <= 65040;
end
1721:begin
x_i <= 65135;
end
1722:begin
x_i <= 65269;
end
1723:begin
x_i <= 65414;
end
1724:begin
x_i <= 20;
end
1725:begin
x_i <= 65476;
end
1726:begin
x_i <= 65224;
end
1727:begin
x_i <= 65057;
end
1728:begin
x_i <= 64943;
end
1729:begin
x_i <= 64876;
end
1730:begin
x_i <= 64731;
end
1731:begin
x_i <= 64824;
end
1732:begin
x_i <= 65141;
end
1733:begin
x_i <= 65475;
end
1734:begin
x_i <= 226;
end
1735:begin
x_i <= 337;
end
1736:begin
x_i <= 382;
end
1737:begin
x_i <= 299;
end
1738:begin
x_i <= 30;
end
1739:begin
x_i <= 65486;
end
1740:begin
x_i <= 65328;
end
1741:begin
x_i <= 65219;
end
1742:begin
x_i <= 65304;
end
1743:begin
x_i <= 65370;
end
1744:begin
x_i <= 65513;
end
1745:begin
x_i <= 88;
end
1746:begin
x_i <= 144;
end
1747:begin
x_i <= 179;
end
1748:begin
x_i <= 101;
end
1749:begin
x_i <= 37;
end
1750:begin
x_i <= 62;
end
1751:begin
x_i <= 96;
end
1752:begin
x_i <= 86;
end
1753:begin
x_i <= 136;
end
1754:begin
x_i <= 295;
end
1755:begin
x_i <= 450;
end
1756:begin
x_i <= 484;
end
1757:begin
x_i <= 490;
end
1758:begin
x_i <= 527;
end
1759:begin
x_i <= 417;
end
1760:begin
x_i <= 416;
end
1761:begin
x_i <= 458;
end
1762:begin
x_i <= 611;
end
1763:begin
x_i <= 793;
end
1764:begin
x_i <= 346;
end
1765:begin
x_i <= 65125;
end
1766:begin
x_i <= 64834;
end
1767:begin
x_i <= 64995;
end
1768:begin
x_i <= 65264;
end
1769:begin
x_i <= 65491;
end
1770:begin
x_i <= 159;
end
1771:begin
x_i <= 490;
end
1772:begin
x_i <= 211;
end
1773:begin
x_i <= 65324;
end
1774:begin
x_i <= 65458;
end
1775:begin
x_i <= 65399;
end
1776:begin
x_i <= 65017;
end
1777:begin
x_i <= 64811;
end
1778:begin
x_i <= 65009;
end
1779:begin
x_i <= 65310;
end
1780:begin
x_i <= 65411;
end
1781:begin
x_i <= 210;
end
1782:begin
x_i <= 658;
end
1783:begin
x_i <= 486;
end
1784:begin
x_i <= 160;
end
1785:begin
x_i <= 79;
end
1786:begin
x_i <= 35;
end
1787:begin
x_i <= 65363;
end
1788:begin
x_i <= 65248;
end
1789:begin
x_i <= 65327;
end
1790:begin
x_i <= 65454;
end
1791:begin
x_i <= 65435;
end
1792:begin
x_i <= 65470;
end
1793:begin
x_i <= 88;
end
1794:begin
x_i <= 65412;
end
1795:begin
x_i <= 64961;
end
1796:begin
x_i <= 64856;
end
1797:begin
x_i <= 64832;
end
1798:begin
x_i <= 64891;
end
1799:begin
x_i <= 64965;
end
1800:begin
x_i <= 65112;
end
1801:begin
x_i <= 65425;
end
1802:begin
x_i <= 65529;
end
1803:begin
x_i <= 85;
end
1804:begin
x_i <= 227;
end
1805:begin
x_i <= 169;
end
1806:begin
x_i <= 53;
end
1807:begin
x_i <= 65400;
end
1808:begin
x_i <= 65280;
end
1809:begin
x_i <= 65352;
end
1810:begin
x_i <= 65416;
end
1811:begin
x_i <= 65518;
end
1812:begin
x_i <= 88;
end
1813:begin
x_i <= 117;
end
1814:begin
x_i <= 83;
end
1815:begin
x_i <= 68;
end
1816:begin
x_i <= 69;
end
1817:begin
x_i <= 70;
end
1818:begin
x_i <= 34;
end
1819:begin
x_i <= 32;
end
1820:begin
x_i <= 96;
end
1821:begin
x_i <= 177;
end
1822:begin
x_i <= 249;
end
1823:begin
x_i <= 299;
end
1824:begin
x_i <= 346;
end
1825:begin
x_i <= 344;
end
1826:begin
x_i <= 223;
end
1827:begin
x_i <= 203;
end
1828:begin
x_i <= 240;
end
1829:begin
x_i <= 276;
end
1830:begin
x_i <= 292;
end
1831:begin
x_i <= 365;
end
1832:begin
x_i <= 504;
end
1833:begin
x_i <= 658;
end
1834:begin
x_i <= 491;
end
1835:begin
x_i <= 128;
end
1836:begin
x_i <= 65363;
end
1837:begin
x_i <= 65241;
end
1838:begin
x_i <= 65275;
end
1839:begin
x_i <= 65343;
end
1840:begin
x_i <= 65482;
end
1841:begin
x_i <= 147;
end
1842:begin
x_i <= 66;
end
1843:begin
x_i <= 65335;
end
1844:begin
x_i <= 65331;
end
1845:begin
x_i <= 65394;
end
1846:begin
x_i <= 65215;
end
1847:begin
x_i <= 65123;
end
1848:begin
x_i <= 65149;
end
1849:begin
x_i <= 65231;
end
1850:begin
x_i <= 65340;
end
1851:begin
x_i <= 65523;
end
1852:begin
x_i <= 176;
end
1853:begin
x_i <= 189;
end
1854:begin
x_i <= 70;
end
1855:begin
x_i <= 19;
end
1856:begin
x_i <= 65514;
end
1857:begin
x_i <= 65439;
end
1858:begin
x_i <= 65408;
end
1859:begin
x_i <= 65363;
end
1860:begin
x_i <= 65398;
end
1861:begin
x_i <= 65461;
end
1862:begin
x_i <= 42;
end
1863:begin
x_i <= 111;
end
1864:begin
x_i <= 65443;
end
1865:begin
x_i <= 65240;
end
1866:begin
x_i <= 65153;
end
1867:begin
x_i <= 65077;
end
1868:begin
x_i <= 65088;
end
1869:begin
x_i <= 65127;
end
1870:begin
x_i <= 65179;
end
1871:begin
x_i <= 65268;
end
1872:begin
x_i <= 65338;
end
1873:begin
x_i <= 5;
end
1874:begin
x_i <= 156;
end
1875:begin
x_i <= 98;
end
1876:begin
x_i <= 65505;
end
1877:begin
x_i <= 65415;
end
1878:begin
x_i <= 65412;
end
1879:begin
x_i <= 65390;
end
1880:begin
x_i <= 65430;
end
1881:begin
x_i <= 3;
end
1882:begin
x_i <= 26;
end
1883:begin
x_i <= 65;
end
1884:begin
x_i <= 94;
end
1885:begin
x_i <= 171;
end
1886:begin
x_i <= 180;
end
1887:begin
x_i <= 99;
end
1888:begin
x_i <= 14;
end
1889:begin
x_i <= 54;
end
1890:begin
x_i <= 75;
end
1891:begin
x_i <= 109;
end
1892:begin
x_i <= 140;
end
1893:begin
x_i <= 164;
end
1894:begin
x_i <= 135;
end
1895:begin
x_i <= 69;
end
1896:begin
x_i <= 54;
end
1897:begin
x_i <= 52;
end
1898:begin
x_i <= 63;
end
1899:begin
x_i <= 14;
end
1900:begin
x_i <= 21;
end
1901:begin
x_i <= 93;
end
1902:begin
x_i <= 169;
end
1903:begin
x_i <= 216;
end
1904:begin
x_i <= 223;
end
1905:begin
x_i <= 273;
end
1906:begin
x_i <= 291;
end
1907:begin
x_i <= 334;
end
1908:begin
x_i <= 351;
end
1909:begin
x_i <= 213;
end
1910:begin
x_i <= 28;
end
1911:begin
x_i <= 65410;
end
1912:begin
x_i <= 65375;
end
1913:begin
x_i <= 65396;
end
1914:begin
x_i <= 65510;
end
1915:begin
x_i <= 98;
end
1916:begin
x_i <= 68;
end
1917:begin
x_i <= 65476;
end
1918:begin
x_i <= 65471;
end
1919:begin
x_i <= 65449;
end
1920:begin
x_i <= 65332;
end
1921:begin
x_i <= 65284;
end
1922:begin
x_i <= 65299;
end
1923:begin
x_i <= 65318;
end
1924:begin
x_i <= 65316;
end
1925:begin
x_i <= 65476;
end
1926:begin
x_i <= 56;
end
1927:begin
x_i <= 13;
end
1928:begin
x_i <= 65512;
end
1929:begin
x_i <= 65469;
end
1930:begin
x_i <= 65413;
end
1931:begin
x_i <= 65366;
end
1932:begin
x_i <= 65332;
end
1933:begin
x_i <= 65339;
end
1934:begin
x_i <= 65342;
end
1935:begin
x_i <= 65451;
end
1936:begin
x_i <= 65527;
end
1937:begin
x_i <= 52;
end
1938:begin
x_i <= 53;
end
1939:begin
x_i <= 65506;
end
1940:begin
x_i <= 65428;
end
1941:begin
x_i <= 65381;
end
1942:begin
x_i <= 65382;
end
1943:begin
x_i <= 65370;
end
1944:begin
x_i <= 65392;
end
1945:begin
x_i <= 65471;
end
1946:begin
x_i <= 65518;
end
1947:begin
x_i <= 44;
end
1948:begin
x_i <= 83;
end
1949:begin
x_i <= 36;
end
1950:begin
x_i <= 65519;
end
1951:begin
x_i <= 65435;
end
1952:begin
x_i <= 65363;
end
1953:begin
x_i <= 65446;
end
1954:begin
x_i <= 65496;
end
1955:begin
x_i <= 25;
end
1956:begin
x_i <= 62;
end
1957:begin
x_i <= 108;
end
1958:begin
x_i <= 143;
end
1959:begin
x_i <= 124;
end
1960:begin
x_i <= 76;
end
1961:begin
x_i <= 4;
end
1962:begin
x_i <= 65472;
end
1963:begin
x_i <= 65431;
end
1964:begin
x_i <= 65459;
end
1965:begin
x_i <= 65479;
end
1966:begin
x_i <= 65534;
end
1967:begin
x_i <= 80;
end
1968:begin
x_i <= 89;
end
1969:begin
x_i <= 77;
end
1970:begin
x_i <= 40;
end
1971:begin
x_i <= 65509;
end
1972:begin
x_i <= 65428;
end
1973:begin
x_i <= 65379;
end
1974:begin
x_i <= 65439;
end
1975:begin
x_i <= 65464;
end
1976:begin
x_i <= 65534;
end
1977:begin
x_i <= 78;
end
1978:begin
x_i <= 87;
end
1979:begin
x_i <= 41;
end
1980:begin
x_i <= 11;
end
1981:begin
x_i <= 65530;
end
1982:begin
x_i <= 65521;
end
1983:begin
x_i <= 65480;
end
1984:begin
x_i <= 65488;
end
1985:begin
x_i <= 65503;
end
1986:begin
x_i <= 34;
end
1987:begin
x_i <= 74;
end
1988:begin
x_i <= 118;
end
1989:begin
x_i <= 114;
end
1990:begin
x_i <= 160;
end
1991:begin
x_i <= 94;
end
1992:begin
x_i <= 8;
end
1993:begin
x_i <= 65515;
end
1994:begin
x_i <= 65529;
end
1995:begin
x_i <= 65515;
end
1996:begin
x_i <= 65522;
end
1997:begin
x_i <= 30;
end
1998:begin
x_i <= 41;
end
1999:begin
x_i <= 53;
end
2000:begin
x_i <= 58;
end
2001:begin
x_i <= 65512;
end
2002:begin
x_i <= 65474;
end
2003:begin
x_i <= 65429;
end
2004:begin
x_i <= 65368;
end
2005:begin
x_i <= 65400;
end
2006:begin
x_i <= 65425;
end
2007:begin
x_i <= 65452;
end
2008:begin
x_i <= 65472;
end
2009:begin
x_i <= 65506;
end
2010:begin
x_i <= 17;
end
2011:begin
x_i <= 1;
end
2012:begin
x_i <= 65482;
end
2013:begin
x_i <= 65524;
end
2014:begin
x_i <= 65509;
end
2015:begin
x_i <= 65436;
end
2016:begin
x_i <= 65495;
end
2017:begin
x_i <= 65522;
end
2018:begin
x_i <= 65514;
end
2019:begin
x_i <= 65456;
end
2020:begin
x_i <= 65414;
end
2021:begin
x_i <= 65445;
end
2022:begin
x_i <= 65439;
end
2023:begin
x_i <= 65507;
end
2024:begin
x_i <= 65493;
end
2025:begin
x_i <= 65433;
end
2026:begin
x_i <= 65418;
end
2027:begin
x_i <= 65449;
end
2028:begin
x_i <= 65438;
end
2029:begin
x_i <= 65420;
end
2030:begin
x_i <= 65440;
end
2031:begin
x_i <= 65402;
end
2032:begin
x_i <= 65426;
end
2033:begin
x_i <= 65484;
end
2034:begin
x_i <= 65511;
end
2035:begin
x_i <= 8;
end
2036:begin
x_i <= 25;
end
2037:begin
x_i <= 18;
end
2038:begin
x_i <= 65535;
end
2039:begin
x_i <= 65443;
end
2040:begin
x_i <= 65386;
end
2041:begin
x_i <= 65424;
end
2042:begin
x_i <= 65437;
end
2043:begin
x_i <= 65471;
end
2044:begin
x_i <= 65510;
end
2045:begin
x_i <= 36;
end
2046:begin
x_i <= 65529;
end
2047:begin
x_i <= 65491;
end
2048:begin
x_i <= 65470;
end
2049:begin
x_i <= 65418;
end
2050:begin
x_i <= 65422;
end
2051:begin
x_i <= 65431;
end
2052:begin
x_i <= 65474;
end
2053:begin
x_i <= 65485;
end
2054:begin
x_i <= 65513;
end
2055:begin
x_i <= 65532;
end
2056:begin
x_i <= 65533;
end
2057:begin
x_i <= 35;
end
2058:begin
x_i <= 65533;
end
2059:begin
x_i <= 65503;
end
2060:begin
x_i <= 65452;
end
2061:begin
x_i <= 65449;
end
2062:begin
x_i <= 65464;
end
2063:begin
x_i <= 65514;
end
2064:begin
x_i <= 65523;
end
2065:begin
x_i <= 67;
end
2066:begin
x_i <= 41;
end
2067:begin
x_i <= 24;
end
2068:begin
x_i <= 23;
end
2069:begin
x_i <= 56;
end
2070:begin
x_i <= 12;
end
2071:begin
x_i <= 65533;
end
2072:begin
x_i <= 65521;
end
2073:begin
x_i <= 65528;
end
2074:begin
x_i <= 64;
end
2075:begin
x_i <= 67;
end
2076:begin
x_i <= 88;
end
2077:begin
x_i <= 87;
end
2078:begin
x_i <= 36;
end
2079:begin
x_i <= 25;
end
2080:begin
x_i <= 65505;
end
2081:begin
x_i <= 55;
end
2082:begin
x_i <= 42;
end
2083:begin
x_i <= 56;
end
2084:begin
x_i <= 57;
end
2085:begin
x_i <= 64;
end
2086:begin
x_i <= 81;
end
2087:begin
x_i <= 38;
end
2088:begin
x_i <= 65535;
end
2089:begin
x_i <= 65524;
end
2090:begin
x_i <= 65531;
end
2091:begin
x_i <= 65519;
end
2092:begin
x_i <= 4;
end
2093:begin
x_i <= 33;
end
2094:begin
x_i <= 23;
end
2095:begin
x_i <= 65528;
end
2096:begin
x_i <= 65518;
end
2097:begin
x_i <= 65484;
end
2098:begin
x_i <= 65469;
end
2099:begin
x_i <= 65388;
end
2100:begin
x_i <= 65346;
end
2101:begin
x_i <= 65385;
end
2102:begin
x_i <= 65435;
end
2103:begin
x_i <= 65505;
end
2104:begin
x_i <= 65518;
end
2105:begin
x_i <= 22;
end
2106:begin
x_i <= 13;
end
2107:begin
x_i <= 65512;
end
2108:begin
x_i <= 65448;
end
2109:begin
x_i <= 65410;
end
2110:begin
x_i <= 65395;
end
2111:begin
x_i <= 65405;
end
2112:begin
x_i <= 65430;
end
2113:begin
x_i <= 65476;
end
2114:begin
x_i <= 65513;
end
2115:begin
x_i <= 65523;
end
2116:begin
x_i <= 65508;
end
2117:begin
x_i <= 65444;
end
2118:begin
x_i <= 65444;
end
2119:begin
x_i <= 65420;
end
2120:begin
x_i <= 65432;
end
2121:begin
x_i <= 65435;
end
2122:begin
x_i <= 65437;
end
2123:begin
x_i <= 65501;
end
2124:begin
x_i <= 65489;
end
2125:begin
x_i <= 65493;
end
2126:begin
x_i <= 65516;
end
2127:begin
x_i <= 65499;
end
2128:begin
x_i <= 65497;
end
2129:begin
x_i <= 65455;
end
2130:begin
x_i <= 65442;
end
2131:begin
x_i <= 65439;
end
2132:begin
x_i <= 65437;
end
2133:begin
x_i <= 65464;
end
2134:begin
x_i <= 65530;
end
2135:begin
x_i <= 33;
end
2136:begin
x_i <= 43;
end
2137:begin
x_i <= 70;
end
2138:begin
x_i <= 55;
end
2139:begin
x_i <= 65534;
end
2140:begin
x_i <= 65476;
end
2141:begin
x_i <= 65495;
end
2142:begin
x_i <= 65475;
end
2143:begin
x_i <= 65502;
end
2144:begin
x_i <= 8;
end
2145:begin
x_i <= 59;
end
2146:begin
x_i <= 76;
end
2147:begin
x_i <= 72;
end
2148:begin
x_i <= 63;
end
2149:begin
x_i <= 51;
end
2150:begin
x_i <= 22;
end
2151:begin
x_i <= 41;
end
2152:begin
x_i <= 35;
end
2153:begin
x_i <= 30;
end
2154:begin
x_i <= 23;
end
2155:begin
x_i <= 20;
end
2156:begin
x_i <= 22;
end
2157:begin
x_i <= 56;
end
2158:begin
x_i <= 54;
end
2159:begin
x_i <= 51;
end
2160:begin
x_i <= 40;
end
2161:begin
x_i <= 32;
end
2162:begin
x_i <= 34;
end
2163:begin
x_i <= 9;
end
2164:begin
x_i <= 65520;
end
2165:begin
x_i <= 65520;
end
2166:begin
x_i <= 65485;
end
2167:begin
x_i <= 65460;
end
2168:begin
x_i <= 65464;
end
2169:begin
x_i <= 65456;
end
2170:begin
x_i <= 65508;
end
2171:begin
x_i <= 65517;
end
2172:begin
x_i <= 65533;
end
2173:begin
x_i <= 65519;
end
2174:begin
x_i <= 65517;
end
2175:begin
x_i <= 65532;
end
2176:begin
x_i <= 65480;
end
2177:begin
x_i <= 65446;
end
2178:begin
x_i <= 65418;
end
2179:begin
x_i <= 65459;
end
2180:begin
x_i <= 65447;
end
2181:begin
x_i <= 65487;
end
2182:begin
x_i <= 65523;
end
2183:begin
x_i <= 11;
end
2184:begin
x_i <= 0;
end
2185:begin
x_i <= 65514;
end
2186:begin
x_i <= 65511;
end
2187:begin
x_i <= 65470;
end
2188:begin
x_i <= 65462;
end
2189:begin
x_i <= 65450;
end
2190:begin
x_i <= 65469;
end
2191:begin
x_i <= 65483;
end
2192:begin
x_i <= 65525;
end
2193:begin
x_i <= 23;
end
2194:begin
x_i <= 65534;
end
2195:begin
x_i <= 65525;
end
2196:begin
x_i <= 65499;
end
2197:begin
x_i <= 65509;
end
2198:begin
x_i <= 65478;
end
2199:begin
x_i <= 65460;
end
2200:begin
x_i <= 65466;
end
2201:begin
x_i <= 65442;
end
2202:begin
x_i <= 65471;
end
2203:begin
x_i <= 65515;
end
2204:begin
x_i <= 14;
end
2205:begin
x_i <= 21;
end
2206:begin
x_i <= 14;
end
2207:begin
x_i <= 65533;
end
2208:begin
x_i <= 65495;
end
2209:begin
x_i <= 10;
end
2210:begin
x_i <= 65481;
end
2211:begin
x_i <= 65489;
end
2212:begin
x_i <= 65500;
end
2213:begin
x_i <= 65517;
end
2214:begin
x_i <= 18;
end
2215:begin
x_i <= 24;
end
2216:begin
x_i <= 63;
end
2217:begin
x_i <= 62;
end
2218:begin
x_i <= 66;
end
2219:begin
x_i <= 49;
end
2220:begin
x_i <= 49;
end
2221:begin
x_i <= 66;
end
2222:begin
x_i <= 26;
end
2223:begin
x_i <= 65523;
end
2224:begin
x_i <= 65526;
end
2225:begin
x_i <= 65489;
end
2226:begin
x_i <= 65521;
end
2227:begin
x_i <= 10;
end
2228:begin
x_i <= 15;
end
2229:begin
x_i <= 34;
end
2230:begin
x_i <= 48;
end
2231:begin
x_i <= 55;
end
2232:begin
x_i <= 28;
end
2233:begin
x_i <= 8;
end
2234:begin
x_i <= 65533;
end
2235:begin
x_i <= 65474;
end
2236:begin
x_i <= 65432;
end
2237:begin
x_i <= 65466;
end
2238:begin
x_i <= 65441;
end
2239:begin
x_i <= 65513;
end
2240:begin
x_i <= 65508;
end
2241:begin
x_i <= 65513;
end
2242:begin
x_i <= 65512;
end
2243:begin
x_i <= 65510;
end
2244:begin
x_i <= 65506;
end
2245:begin
x_i <= 65480;
end
2246:begin
x_i <= 65483;
end
2247:begin
x_i <= 65438;
end
2248:begin
x_i <= 65418;
end
2249:begin
x_i <= 65466;
end
2250:begin
x_i <= 65493;
end
2251:begin
x_i <= 65510;
end
2252:begin
x_i <= 65524;
end
2253:begin
x_i <= 65524;
end
2254:begin
x_i <= 65499;
end
2255:begin
x_i <= 65489;
end
2256:begin
x_i <= 65495;
end
2257:begin
x_i <= 65458;
end
2258:begin
x_i <= 65479;
end
2259:begin
x_i <= 65478;
end
2260:begin
x_i <= 65472;
end
2261:begin
x_i <= 65513;
end
2262:begin
x_i <= 65519;
end
2263:begin
x_i <= 65535;
end
2264:begin
x_i <= 65521;
end
2265:begin
x_i <= 65527;
end
2266:begin
x_i <= 5;
end
2267:begin
x_i <= 65503;
end
2268:begin
x_i <= 65496;
end
2269:begin
x_i <= 65483;
end
2270:begin
x_i <= 65470;
end
2271:begin
x_i <= 65473;
end
2272:begin
x_i <= 65505;
end
2273:begin
x_i <= 0;
end
2274:begin
x_i <= 65534;
end
2275:begin
x_i <= 18;
end
2276:begin
x_i <= 65528;
end
2277:begin
x_i <= 0;
end
2278:begin
x_i <= 12;
end
2279:begin
x_i <= 6;
end
2280:begin
x_i <= 65511;
end
2281:begin
x_i <= 65518;
end
2282:begin
x_i <= 3;
end
2283:begin
x_i <= 65525;
end
2284:begin
x_i <= 17;
end
2285:begin
x_i <= 41;
end
2286:begin
x_i <= 70;
end
2287:begin
x_i <= 45;
end
2288:begin
x_i <= 61;
end
2289:begin
x_i <= 19;
end
2290:begin
x_i <= 18;
end
2291:begin
x_i <= 65522;
end
2292:begin
x_i <= 3;
end
2293:begin
x_i <= 65516;
end
2294:begin
x_i <= 65507;
end
2295:begin
x_i <= 65532;
end
2296:begin
x_i <= 65526;
end
2297:begin
x_i <= 65517;
end
2298:begin
x_i <= 65524;
end
2299:begin
x_i <= 65492;
end
2300:begin
x_i <= 65496;
end
2301:begin
x_i <= 65490;
end
2302:begin
x_i <= 65439;
end
2303:begin
x_i <= 65459;
end
2304:begin
x_i <= 65482;
end
2305:begin
x_i <= 65501;
end
2306:begin
x_i <= 65483;
end
2307:begin
x_i <= 65497;
end
2308:begin
x_i <= 65530;
end
2309:begin
x_i <= 65493;
end
2310:begin
x_i <= 65461;
end
2311:begin
x_i <= 65481;
end
2312:begin
x_i <= 65479;
end
2313:begin
x_i <= 65480;
end
2314:begin
x_i <= 65462;
end
2315:begin
x_i <= 65495;
end
2316:begin
x_i <= 65498;
end
2317:begin
x_i <= 65501;
end
2318:begin
x_i <= 65479;
end
2319:begin
x_i <= 65495;
end
2320:begin
x_i <= 65496;
end
2321:begin
x_i <= 65491;
end
2322:begin
x_i <= 65473;
end
2323:begin
x_i <= 65497;
end
2324:begin
x_i <= 65481;
end
2325:begin
x_i <= 65498;
end
2326:begin
x_i <= 65505;
end
2327:begin
x_i <= 41;
end
2328:begin
x_i <= 39;
end
2329:begin
x_i <= 21;
end
2330:begin
x_i <= 7;
end
2331:begin
x_i <= 3;
end
2332:begin
x_i <= 65512;
end
2333:begin
x_i <= 65462;
end
2334:begin
x_i <= 65481;
end
2335:begin
x_i <= 65483;
end
2336:begin
x_i <= 65487;
end
2337:begin
x_i <= 65450;
end
2338:begin
x_i <= 65514;
end
2339:begin
x_i <= 65502;
end
2340:begin
x_i <= 65514;
end
2341:begin
x_i <= 27;
end
2342:begin
x_i <= 18;
end
2343:begin
x_i <= 65518;
end
2344:begin
x_i <= 65522;
end
2345:begin
x_i <= 65515;
end
2346:begin
x_i <= 65477;
end
2347:begin
x_i <= 65500;
end
2348:begin
x_i <= 65496;
end
2349:begin
x_i <= 65518;
end
2350:begin
x_i <= 65509;
end
2351:begin
x_i <= 65518;
end
2352:begin
x_i <= 3;
end
2353:begin
x_i <= 65529;
end
2354:begin
x_i <= 65517;
end
2355:begin
x_i <= 23;
end
2356:begin
x_i <= 17;
end
2357:begin
x_i <= 29;
end
2358:begin
x_i <= 25;
end
2359:begin
x_i <= 65526;
end
2360:begin
x_i <= 65525;
end
2361:begin
x_i <= 65520;
end
2362:begin
x_i <= 65513;
end
2363:begin
x_i <= 65535;
end
2364:begin
x_i <= 5;
end
2365:begin
x_i <= 19;
end
2366:begin
x_i <= 65521;
end
2367:begin
x_i <= 65511;
end
2368:begin
x_i <= 65491;
end
2369:begin
x_i <= 65482;
end
2370:begin
x_i <= 65475;
end
2371:begin
x_i <= 65457;
end
2372:begin
x_i <= 65465;
end
2373:begin
x_i <= 65464;
end
2374:begin
x_i <= 65472;
end
2375:begin
x_i <= 65492;
end
2376:begin
x_i <= 65529;
end
2377:begin
x_i <= 65506;
end
2378:begin
x_i <= 9;
end
2379:begin
x_i <= 65500;
end
2380:begin
x_i <= 65490;
end
2381:begin
x_i <= 65495;
end
2382:begin
x_i <= 65460;
end
2383:begin
x_i <= 65472;
end
2384:begin
x_i <= 65496;
end
2385:begin
x_i <= 65466;
end
2386:begin
x_i <= 65475;
end
2387:begin
x_i <= 65499;
end
2388:begin
x_i <= 0;
end
2389:begin
x_i <= 65490;
end
2390:begin
x_i <= 65520;
end
2391:begin
x_i <= 65462;
end
2392:begin
x_i <= 65455;
end
2393:begin
x_i <= 65441;
end
2394:begin
x_i <= 65448;
end
2395:begin
x_i <= 65487;
end
2396:begin
x_i <= 65511;
end
2397:begin
x_i <= 65513;
end
2398:begin
x_i <= 13;
end
2399:begin
x_i <= 6;
end
2400:begin
x_i <= 65528;
end
2401:begin
x_i <= 65495;
end
2402:begin
x_i <= 65496;
end
2403:begin
x_i <= 65431;
end
2404:begin
x_i <= 65441;
end
2405:begin
x_i <= 65471;
end
2406:begin
x_i <= 65477;
end
2407:begin
x_i <= 65469;
end
2408:begin
x_i <= 65496;
end
2409:begin
x_i <= 65459;
end
2410:begin
x_i <= 65497;
end
2411:begin
x_i <= 65525;
end
2412:begin
x_i <= 65531;
end
2413:begin
x_i <= 65524;
end
2414:begin
x_i <= 65534;
end
2415:begin
x_i <= 65515;
end
2416:begin
x_i <= 65499;
end
2417:begin
x_i <= 65504;
end
2418:begin
x_i <= 65506;
end
2419:begin
x_i <= 19;
end
2420:begin
x_i <= 8;
end
2421:begin
x_i <= 6;
end
2422:begin
x_i <= 65534;
end
2423:begin
x_i <= 65535;
end
2424:begin
x_i <= 65522;
end
2425:begin
x_i <= 21;
end
2426:begin
x_i <= 65473;
end
2427:begin
x_i <= 65512;
end
2428:begin
x_i <= 65523;
end
2429:begin
x_i <= 65519;
end
2430:begin
x_i <= 65528;
end
2431:begin
x_i <= 65525;
end
2432:begin
x_i <= 36;
end
2433:begin
x_i <= 11;
end
2434:begin
x_i <= 2;
end
2435:begin
x_i <= 16;
end
2436:begin
x_i <= 3;
end
2437:begin
x_i <= 65493;
end
2438:begin
x_i <= 65451;
end
2439:begin
x_i <= 65483;
end
2440:begin
x_i <= 65508;
end
2441:begin
x_i <= 65515;
end
2442:begin
x_i <= 65487;
end
2443:begin
x_i <= 65484;
end
2444:begin
x_i <= 65506;
end
2445:begin
x_i <= 65505;
end
2446:begin
x_i <= 5;
end
2447:begin
x_i <= 1;
end
2448:begin
x_i <= 5;
end
2449:begin
x_i <= 65502;
end
2450:begin
x_i <= 65517;
end
2451:begin
x_i <= 65509;
end
2452:begin
x_i <= 65519;
end
2453:begin
x_i <= 19;
end
2454:begin
x_i <= 65521;
end
2455:begin
x_i <= 26;
end
2456:begin
x_i <= 65526;
end
2457:begin
x_i <= 65517;
end
2458:begin
x_i <= 65506;
end
2459:begin
x_i <= 65525;
end
2460:begin
x_i <= 65487;
end
2461:begin
x_i <= 65457;
end
2462:begin
x_i <= 65445;
end
2463:begin
x_i <= 65453;
end
2464:begin
x_i <= 65499;
end
2465:begin
x_i <= 65494;
end
2466:begin
x_i <= 65513;
end
2467:begin
x_i <= 65508;
end
2468:begin
x_i <= 65511;
end
2469:begin
x_i <= 16;
end
2470:begin
x_i <= 7;
end
2471:begin
x_i <= 65519;
end
2472:begin
x_i <= 65458;
end
2473:begin
x_i <= 65444;
end
2474:begin
x_i <= 65448;
end
2475:begin
x_i <= 65463;
end
2476:begin
x_i <= 65463;
end
2477:begin
x_i <= 65459;
end
2478:begin
x_i <= 65465;
end
2479:begin
x_i <= 65473;
end
2480:begin
x_i <= 65481;
end
2481:begin
x_i <= 65487;
end
2482:begin
x_i <= 65516;
end
2483:begin
x_i <= 65516;
end
2484:begin
x_i <= 65505;
end
2485:begin
x_i <= 65505;
end
2486:begin
x_i <= 65527;
end
2487:begin
x_i <= 65501;
end
2488:begin
x_i <= 65532;
end
2489:begin
x_i <= 65532;
end
2490:begin
x_i <= 65530;
end
2491:begin
x_i <= 65522;
end
2492:begin
x_i <= 65496;
end
2493:begin
x_i <= 65532;
end
2494:begin
x_i <= 65478;
end
2495:begin
x_i <= 65493;
end
2496:begin
x_i <= 65463;
end
2497:begin
x_i <= 65495;
end
2498:begin
x_i <= 65488;
end
2499:begin
x_i <= 65513;
end
2500:begin
x_i <= 18;
end
2501:begin
x_i <= 24;
end
2502:begin
x_i <= 29;
end
2503:begin
x_i <= 14;
end
2504:begin
x_i <= 5;
end
2505:begin
x_i <= 65520;
end
2506:begin
x_i <= 65505;
end
2507:begin
x_i <= 65482;
end
2508:begin
x_i <= 65482;
end
2509:begin
x_i <= 65482;
end
2510:begin
x_i <= 65496;
end
2511:begin
x_i <= 65490;
end
2512:begin
x_i <= 65498;
end
2513:begin
x_i <= 65497;
end
2514:begin
x_i <= 65496;
end
2515:begin
x_i <= 65524;
end
2516:begin
x_i <= 65523;
end
2517:begin
x_i <= 65518;
end
2518:begin
x_i <= 65505;
end
2519:begin
x_i <= 65507;
end
2520:begin
x_i <= 65512;
end
2521:begin
x_i <= 65519;
end
2522:begin
x_i <= 65504;
end
2523:begin
x_i <= 65496;
end
2524:begin
x_i <= 4;
end
2525:begin
x_i <= 65507;
end
2526:begin
x_i <= 65498;
end
2527:begin
x_i <= 65533;
end
2528:begin
x_i <= 65476;
end
2529:begin
x_i <= 65470;
end
2530:begin
x_i <= 65512;
end
2531:begin
x_i <= 65496;
end
2532:begin
x_i <= 65509;
end
2533:begin
x_i <= 65515;
end
2534:begin
x_i <= 65504;
end
2535:begin
x_i <= 65495;
end
2536:begin
x_i <= 65512;
end
2537:begin
x_i <= 65506;
end
2538:begin
x_i <= 65505;
end
2539:begin
x_i <= 65515;
end
2540:begin
x_i <= 65510;
end
2541:begin
x_i <= 65494;
end
2542:begin
x_i <= 65495;
end
2543:begin
x_i <= 65485;
end
2544:begin
x_i <= 65484;
end
2545:begin
x_i <= 65498;
end
2546:begin
x_i <= 65486;
end
2547:begin
x_i <= 65489;
end
2548:begin
x_i <= 65462;
end
2549:begin
x_i <= 65462;
end
2550:begin
x_i <= 65503;
end
2551:begin
x_i <= 65500;
end
2552:begin
x_i <= 65500;
end
2553:begin
x_i <= 65508;
end
2554:begin
x_i <= 65506;
end
2555:begin
x_i <= 65517;
end
2556:begin
x_i <= 65500;
end
2557:begin
x_i <= 65520;
end
2558:begin
x_i <= 65513;
end
2559:begin
x_i <= 65532;
end
2560:begin
x_i <= 65507;
end
2561:begin
x_i <= 65519;
end
2562:begin
x_i <= 65522;
end
2563:begin
x_i <= 65515;
end
2564:begin
x_i <= 65489;
end
2565:begin
x_i <= 65475;
end
2566:begin
x_i <= 65478;
end
2567:begin
x_i <= 65483;
end
2568:begin
x_i <= 65510;
end
2569:begin
x_i <= 65535;
end
2570:begin
x_i <= 65478;
end
2571:begin
x_i <= 65498;
end
2572:begin
x_i <= 4;
end
2573:begin
x_i <= 38;
end
2574:begin
x_i <= 13;
end
2575:begin
x_i <= 1;
end
2576:begin
x_i <= 65527;
end
2577:begin
x_i <= 65521;
end
2578:begin
x_i <= 65516;
end
2579:begin
x_i <= 65528;
end
2580:begin
x_i <= 65501;
end
2581:begin
x_i <= 65504;
end
2582:begin
x_i <= 65478;
end
2583:begin
x_i <= 65464;
end
2584:begin
x_i <= 65490;
end
2585:begin
x_i <= 65530;
end
2586:begin
x_i <= 65513;
end
2587:begin
x_i <= 65503;
end
2588:begin
x_i <= 65502;
end
2589:begin
x_i <= 65500;
end
2590:begin
x_i <= 65531;
end
2591:begin
x_i <= 2;
end
2592:begin
x_i <= 65513;
end
2593:begin
x_i <= 65500;
end
2594:begin
x_i <= 65505;
end
2595:begin
x_i <= 65516;
end
2596:begin
x_i <= 65479;
end
2597:begin
x_i <= 65477;
end
2598:begin
x_i <= 65482;
end
2599:begin
x_i <= 65494;
end
2600:begin
x_i <= 65494;
end
2601:begin
x_i <= 65507;
end
2602:begin
x_i <= 65498;
end
2603:begin
x_i <= 65522;
end
2604:begin
x_i <= 65495;
end
2605:begin
x_i <= 65494;
end
2606:begin
x_i <= 65481;
end
2607:begin
x_i <= 65487;
end
2608:begin
x_i <= 65475;
end
2609:begin
x_i <= 65486;
end
2610:begin
x_i <= 65489;
end
2611:begin
x_i <= 65523;
end
2612:begin
x_i <= 65504;
end
2613:begin
x_i <= 4;
end
2614:begin
x_i <= 13;
end
2615:begin
x_i <= 65498;
end
2616:begin
x_i <= 65482;
end
2617:begin
x_i <= 65454;
end
2618:begin
x_i <= 65479;
end
2619:begin
x_i <= 65496;
end
2620:begin
x_i <= 65476;
end
2621:begin
x_i <= 65471;
end
2622:begin
x_i <= 65523;
end
2623:begin
x_i <= 65520;
end
2624:begin
x_i <= 65509;
end
2625:begin
x_i <= 65525;
end
2626:begin
x_i <= 6;
end
2627:begin
x_i <= 23;
end
2628:begin
x_i <= 65519;
end
2629:begin
x_i <= 17;
end
2630:begin
x_i <= 4;
end
2631:begin
x_i <= 10;
end
2632:begin
x_i <= 6;
end
2633:begin
x_i <= 65512;
end
2634:begin
x_i <= 65485;
end
2635:begin
x_i <= 65492;
end
2636:begin
x_i <= 65527;
end
2637:begin
x_i <= 65535;
end
2638:begin
x_i <= 0;
end
2639:begin
x_i <= 65528;
end
2640:begin
x_i <= 65525;
end
2641:begin
x_i <= 65529;
end
2642:begin
x_i <= 22;
end
2643:begin
x_i <= 65530;
end
2644:begin
x_i <= 65530;
end
2645:begin
x_i <= 65521;
end
2646:begin
x_i <= 65527;
end
2647:begin
x_i <= 65535;
end
2648:begin
x_i <= 16;
end
2649:begin
x_i <= 20;
end
2650:begin
x_i <= 65535;
end
2651:begin
x_i <= 65517;
end
2652:begin
x_i <= 65505;
end
2653:begin
x_i <= 65519;
end
2654:begin
x_i <= 15;
end
2655:begin
x_i <= 65510;
end
2656:begin
x_i <= 65496;
end
2657:begin
x_i <= 65514;
end
2658:begin
x_i <= 65507;
end
2659:begin
x_i <= 65531;
end
2660:begin
x_i <= 46;
end
2661:begin
x_i <= 12;
end
2662:begin
x_i <= 19;
end
2663:begin
x_i <= 7;
end
2664:begin
x_i <= 65534;
end
2665:begin
x_i <= 65501;
end
2666:begin
x_i <= 65524;
end
2667:begin
x_i <= 65501;
end
2668:begin
x_i <= 65496;
end
2669:begin
x_i <= 65503;
end
2670:begin
x_i <= 65530;
end
2671:begin
x_i <= 18;
end
2672:begin
x_i <= 65527;
end
2673:begin
x_i <= 20;
end
2674:begin
x_i <= 13;
end
2675:begin
x_i <= 65502;
end
2676:begin
x_i <= 65478;
end
2677:begin
x_i <= 65491;
end
2678:begin
x_i <= 65494;
end
2679:begin
x_i <= 65482;
end
2680:begin
x_i <= 65517;
end
2681:begin
x_i <= 65505;
end
2682:begin
x_i <= 65511;
end
2683:begin
x_i <= 65511;
end
2684:begin
x_i <= 65504;
end
2685:begin
x_i <= 65530;
end
2686:begin
x_i <= 65531;
end
2687:begin
x_i <= 65505;
end
2688:begin
x_i <= 65489;
end
2689:begin
x_i <= 65489;
end
2690:begin
x_i <= 65489;
end
2691:begin
x_i <= 65492;
end
2692:begin
x_i <= 65494;
end
2693:begin
x_i <= 65509;
end
2694:begin
x_i <= 65531;
end
2695:begin
x_i <= 65501;
end
2696:begin
x_i <= 65511;
end
2697:begin
x_i <= 65535;
end
2698:begin
x_i <= 3;
end
2699:begin
x_i <= 65519;
end
2700:begin
x_i <= 65528;
end
2701:begin
x_i <= 65519;
end
2702:begin
x_i <= 65473;
end
2703:begin
x_i <= 65473;
end
2704:begin
x_i <= 65486;
end
2705:begin
x_i <= 65489;
end
2706:begin
x_i <= 65500;
end
2707:begin
x_i <= 65487;
end
2708:begin
x_i <= 65514;
end
2709:begin
x_i <= 65524;
end
2710:begin
x_i <= 65505;
end
2711:begin
x_i <= 65532;
end
2712:begin
x_i <= 65522;
end
2713:begin
x_i <= 5;
end
2714:begin
x_i <= 65508;
end
2715:begin
x_i <= 65523;
end
2716:begin
x_i <= 65494;
end
2717:begin
x_i <= 65501;
end
2718:begin
x_i <= 65519;
end
2719:begin
x_i <= 2;
end
2720:begin
x_i <= 65520;
end
2721:begin
x_i <= 65527;
end
2722:begin
x_i <= 65528;
end
2723:begin
x_i <= 65518;
end
2724:begin
x_i <= 65491;
end
2725:begin
x_i <= 65500;
end
2726:begin
x_i <= 65528;
end
2727:begin
x_i <= 65495;
end
2728:begin
x_i <= 65499;
end
2729:begin
x_i <= 65526;
end
2730:begin
x_i <= 65513;
end
2731:begin
x_i <= 19;
end
2732:begin
x_i <= 65534;
end
2733:begin
x_i <= 15;
end
2734:begin
x_i <= 65510;
end
2735:begin
x_i <= 65521;
end
2736:begin
x_i <= 65520;
end
2737:begin
x_i <= 65515;
end
2738:begin
x_i <= 65503;
end
2739:begin
x_i <= 65524;
end
2740:begin
x_i <= 65510;
end
2741:begin
x_i <= 65522;
end
2742:begin
x_i <= 65520;
end
2743:begin
x_i <= 53;
end
2744:begin
x_i <= 4;
end
2745:begin
x_i <= 65522;
end
2746:begin
x_i <= 65524;
end
2747:begin
x_i <= 65489;
end
2748:begin
x_i <= 65493;
end
2749:begin
x_i <= 65489;
end
2750:begin
x_i <= 65507;
end
2751:begin
x_i <= 65512;
end
2752:begin
x_i <= 65492;
end
2753:begin
x_i <= 65509;
end
2754:begin
x_i <= 65530;
end
2755:begin
x_i <= 65521;
end
2756:begin
x_i <= 65513;
end
2757:begin
x_i <= 65502;
end
2758:begin
x_i <= 65488;
end
2759:begin
x_i <= 65481;
end
2760:begin
x_i <= 65498;
end
2761:begin
x_i <= 65461;
end
2762:begin
x_i <= 65484;
end
2763:begin
x_i <= 65501;
end
2764:begin
x_i <= 65518;
end
2765:begin
x_i <= 65506;
end
2766:begin
x_i <= 65524;
end
2767:begin
x_i <= 1;
end
2768:begin
x_i <= 65512;
end
2769:begin
x_i <= 65501;
end
2770:begin
x_i <= 65494;
end
2771:begin
x_i <= 65491;
end
2772:begin
x_i <= 65486;
end
2773:begin
x_i <= 65490;
end
2774:begin
x_i <= 65466;
end
2775:begin
x_i <= 65488;
end
2776:begin
x_i <= 65506;
end
2777:begin
x_i <= 65512;
end
2778:begin
x_i <= 65517;
end
2779:begin
x_i <= 65468;
end
2780:begin
x_i <= 65521;
end
2781:begin
x_i <= 65503;
end
2782:begin
x_i <= 65485;
end
2783:begin
x_i <= 65472;
end
2784:begin
x_i <= 65499;
end
2785:begin
x_i <= 65474;
end
2786:begin
x_i <= 65496;
end
2787:begin
x_i <= 65506;
end
2788:begin
x_i <= 7;
end
2789:begin
x_i <= 65512;
end
2790:begin
x_i <= 0;
end
2791:begin
x_i <= 65518;
end
2792:begin
x_i <= 65497;
end
2793:begin
x_i <= 65492;
end
2794:begin
x_i <= 65457;
end
2795:begin
x_i <= 65453;
end
2796:begin
x_i <= 65491;
end
2797:begin
x_i <= 65494;
end
2798:begin
x_i <= 65524;
end
2799:begin
x_i <= 5;
end
2800:begin
x_i <= 16;
end
2801:begin
x_i <= 65530;
end
2802:begin
x_i <= 65531;
end
2803:begin
x_i <= 65501;
end
2804:begin
x_i <= 65503;
end
2805:begin
x_i <= 65467;
end
2806:begin
x_i <= 65474;
end
2807:begin
x_i <= 65483;
end
2808:begin
x_i <= 65531;
end
2809:begin
x_i <= 65510;
end
2810:begin
x_i <= 11;
end
2811:begin
x_i <= 65516;
end
2812:begin
x_i <= 65506;
end
2813:begin
x_i <= 65502;
end
2814:begin
x_i <= 65496;
end
2815:begin
x_i <= 65475;
end
2816:begin
x_i <= 65470;
end
2817:begin
x_i <= 65490;
end
2818:begin
x_i <= 65492;
end
2819:begin
x_i <= 65491;
end
2820:begin
x_i <= 65486;
end
2821:begin
x_i <= 8;
end
2822:begin
x_i <= 65511;
end
2823:begin
x_i <= 65534;
end
2824:begin
x_i <= 65534;
end
2825:begin
x_i <= 65511;
end
2826:begin
x_i <= 65505;
end
2827:begin
x_i <= 65495;
end
2828:begin
x_i <= 65478;
end
2829:begin
x_i <= 65494;
end
2830:begin
x_i <= 65532;
end
2831:begin
x_i <= 3;
end
2832:begin
x_i <= 15;
end
2833:begin
x_i <= 16;
end
2834:begin
x_i <= 8;
end
2835:begin
x_i <= 26;
end
2836:begin
x_i <= 14;
end
2837:begin
x_i <= 65531;
end
2838:begin
x_i <= 65508;
end
2839:begin
x_i <= 65518;
end
2840:begin
x_i <= 65476;
end
2841:begin
x_i <= 65496;
end
2842:begin
x_i <= 9;
end
2843:begin
x_i <= 113;
end
2844:begin
x_i <= 65481;
end
2845:begin
x_i <= 65284;
end
2846:begin
x_i <= 65360;
end
2847:begin
x_i <= 65400;
end
2848:begin
x_i <= 65405;
end
2849:begin
x_i <= 88;
end
2850:begin
x_i <= 260;
end
2851:begin
x_i <= 225;
end
2852:begin
x_i <= 12;
end
2853:begin
x_i <= 65427;
end
2854:begin
x_i <= 65368;
end
2855:begin
x_i <= 65240;
end
2856:begin
x_i <= 65323;
end
2857:begin
x_i <= 65508;
end
2858:begin
x_i <= 101;
end
2859:begin
x_i <= 159;
end
2860:begin
x_i <= 166;
end
2861:begin
x_i <= 131;
end
2862:begin
x_i <= 17;
end
2863:begin
x_i <= 65476;
end
2864:begin
x_i <= 65382;
end
2865:begin
x_i <= 65358;
end
2866:begin
x_i <= 65428;
end
2867:begin
x_i <= 65520;
end
2868:begin
x_i <= 37;
end
2869:begin
x_i <= 120;
end
2870:begin
x_i <= 6;
end
2871:begin
x_i <= 65363;
end
2872:begin
x_i <= 65267;
end
2873:begin
x_i <= 65286;
end
2874:begin
x_i <= 65365;
end
2875:begin
x_i <= 65424;
end
2876:begin
x_i <= 102;
end
2877:begin
x_i <= 165;
end
2878:begin
x_i <= 102;
end
2879:begin
x_i <= 33;
end
2880:begin
x_i <= 65429;
end
2881:begin
x_i <= 65303;
end
2882:begin
x_i <= 65324;
end
2883:begin
x_i <= 65455;
end
2884:begin
x_i <= 65509;
end
2885:begin
x_i <= 103;
end
2886:begin
x_i <= 198;
end
2887:begin
x_i <= 195;
end
2888:begin
x_i <= 64;
end
2889:begin
x_i <= 12;
end
2890:begin
x_i <= 65482;
end
2891:begin
x_i <= 65452;
end
2892:begin
x_i <= 65497;
end
2893:begin
x_i <= 56;
end
2894:begin
x_i <= 114;
end
2895:begin
x_i <= 155;
end
2896:begin
x_i <= 139;
end
2897:begin
x_i <= 48;
end
2898:begin
x_i <= 7;
end
2899:begin
x_i <= 65457;
end
2900:begin
x_i <= 65445;
end
2901:begin
x_i <= 65421;
end
2902:begin
x_i <= 65528;
end
2903:begin
x_i <= 51;
end
2904:begin
x_i <= 103;
end
2905:begin
x_i <= 145;
end
2906:begin
x_i <= 154;
end
2907:begin
x_i <= 33;
end
2908:begin
x_i <= 65449;
end
2909:begin
x_i <= 65454;
end
2910:begin
x_i <= 65245;
end
2911:begin
x_i <= 65284;
end
2912:begin
x_i <= 65415;
end
2913:begin
x_i <= 65494;
end
2914:begin
x_i <= 65527;
end
2915:begin
x_i <= 82;
end
2916:begin
x_i <= 134;
end
2917:begin
x_i <= 65497;
end
2918:begin
x_i <= 65380;
end
2919:begin
x_i <= 65415;
end
2920:begin
x_i <= 65323;
end
2921:begin
x_i <= 65323;
end
2922:begin
x_i <= 65487;
end
2923:begin
x_i <= 55;
end
2924:begin
x_i <= 20;
end
2925:begin
x_i <= 132;
end
2926:begin
x_i <= 123;
end
2927:begin
x_i <= 65528;
end
2928:begin
x_i <= 65469;
end
2929:begin
x_i <= 65473;
end
2930:begin
x_i <= 65391;
end
2931:begin
x_i <= 65465;
end
2932:begin
x_i <= 28;
end
2933:begin
x_i <= 59;
end
2934:begin
x_i <= 19;
end
2935:begin
x_i <= 65464;
end
2936:begin
x_i <= 65440;
end
2937:begin
x_i <= 65373;
end
2938:begin
x_i <= 65415;
end
2939:begin
x_i <= 65526;
end
2940:begin
x_i <= 176;
end
2941:begin
x_i <= 439;
end
2942:begin
x_i <= 65484;
end
2943:begin
x_i <= 65480;
end
2944:begin
x_i <= 65338;
end
2945:begin
x_i <= 65140;
end
2946:begin
x_i <= 65064;
end
2947:begin
x_i <= 1;
end
2948:begin
x_i <= 232;
end
2949:begin
x_i <= 271;
end
2950:begin
x_i <= 357;
end
2951:begin
x_i <= 246;
end
2952:begin
x_i <= 65439;
end
2953:begin
x_i <= 65087;
end
2954:begin
x_i <= 65123;
end
2955:begin
x_i <= 65051;
end
2956:begin
x_i <= 65300;
end
2957:begin
x_i <= 296;
end
2958:begin
x_i <= 337;
end
2959:begin
x_i <= 316;
end
2960:begin
x_i <= 200;
end
2961:begin
x_i <= 65373;
end
2962:begin
x_i <= 64885;
end
2963:begin
x_i <= 65078;
end
2964:begin
x_i <= 65118;
end
2965:begin
x_i <= 65271;
end
2966:begin
x_i <= 65529;
end
2967:begin
x_i <= 378;
end
2968:begin
x_i <= 288;
end
2969:begin
x_i <= 29;
end
2970:begin
x_i <= 81;
end
2971:begin
x_i <= 65276;
end
2972:begin
x_i <= 65070;
end
2973:begin
x_i <= 65225;
end
2974:begin
x_i <= 65408;
end
2975:begin
x_i <= 65443;
end
2976:begin
x_i <= 203;
end
2977:begin
x_i <= 349;
end
2978:begin
x_i <= 197;
end
2979:begin
x_i <= 106;
end
2980:begin
x_i <= 22;
end
2981:begin
x_i <= 65367;
end
2982:begin
x_i <= 65170;
end
2983:begin
x_i <= 65381;
end
2984:begin
x_i <= 65469;
end
2985:begin
x_i <= 65409;
end
2986:begin
x_i <= 137;
end
2987:begin
x_i <= 129;
end
2988:begin
x_i <= 73;
end
2989:begin
x_i <= 65524;
end
2990:begin
x_i <= 9;
end
2991:begin
x_i <= 65399;
end
2992:begin
x_i <= 65441;
end
2993:begin
x_i <= 65456;
end
2994:begin
x_i <= 65439;
end
2995:begin
x_i <= 65518;
end
2996:begin
x_i <= 70;
end
2997:begin
x_i <= 167;
end
2998:begin
x_i <= 84;
end
2999:begin
x_i <= 179;
end
3000:begin
x_i <= 54;
end
3001:begin
x_i <= 12;
end
3002:begin
x_i <= 61;
end
3003:begin
x_i <= 80;
end
3004:begin
x_i <= 21;
end
3005:begin
x_i <= 65517;
end
3006:begin
x_i <= 97;
end
3007:begin
x_i <= 65529;
end
3008:begin
x_i <= 3;
end
3009:begin
x_i <= 65520;
end
3010:begin
x_i <= 65494;
end
3011:begin
x_i <= 65471;
end
3012:begin
x_i <= 51;
end
3013:begin
x_i <= 11;
end
3014:begin
x_i <= 65357;
end
3015:begin
x_i <= 65380;
end
3016:begin
x_i <= 65281;
end
3017:begin
x_i <= 65314;
end
3018:begin
x_i <= 65378;
end
3019:begin
x_i <= 90;
end
3020:begin
x_i <= 44;
end
3021:begin
x_i <= 91;
end
3022:begin
x_i <= 76;
end
3023:begin
x_i <= 65507;
end
3024:begin
x_i <= 65349;
end
3025:begin
x_i <= 65253;
end
3026:begin
x_i <= 65377;
end
3027:begin
x_i <= 65397;
end
3028:begin
x_i <= 46;
end
3029:begin
x_i <= 214;
end
3030:begin
x_i <= 289;
end
3031:begin
x_i <= 355;
end
3032:begin
x_i <= 155;
end
3033:begin
x_i <= 65514;
end
3034:begin
x_i <= 65342;
end
3035:begin
x_i <= 65199;
end
3036:begin
x_i <= 65313;
end
3037:begin
x_i <= 65510;
end
3038:begin
x_i <= 169;
end
3039:begin
x_i <= 294;
end
3040:begin
x_i <= 293;
end
3041:begin
x_i <= 210;
end
3042:begin
x_i <= 65488;
end
3043:begin
x_i <= 65291;
end
3044:begin
x_i <= 65155;
end
3045:begin
x_i <= 65158;
end
3046:begin
x_i <= 65303;
end
3047:begin
x_i <= 65529;
end
3048:begin
x_i <= 48;
end
3049:begin
x_i <= 135;
end
3050:begin
x_i <= 158;
end
3051:begin
x_i <= 60;
end
3052:begin
x_i <= 65465;
end
3053:begin
x_i <= 65483;
end
3054:begin
x_i <= 65517;
end
3055:begin
x_i <= 65415;
end
3056:begin
x_i <= 65426;
end
3057:begin
x_i <= 29;
end
3058:begin
x_i <= 185;
end
3059:begin
x_i <= 65454;
end
3060:begin
x_i <= 171;
end
3061:begin
x_i <= 77;
end
3062:begin
x_i <= 65427;
end
3063:begin
x_i <= 65436;
end
3064:begin
x_i <= 48;
end
3065:begin
x_i <= 65484;
end
3066:begin
x_i <= 8;
end
3067:begin
x_i <= 193;
end
3068:begin
x_i <= 73;
end
3069:begin
x_i <= 2;
end
3070:begin
x_i <= 65453;
end
3071:begin
x_i <= 65495;
end
3072:begin
x_i <= 65301;
end
3073:begin
x_i <= 65478;
end
3074:begin
x_i <= 120;
end
3075:begin
x_i <= 87;
end
3076:begin
x_i <= 86;
end
3077:begin
x_i <= 177;
end
3078:begin
x_i <= 65368;
end
3079:begin
x_i <= 65138;
end
3080:begin
x_i <= 65282;
end
3081:begin
x_i <= 65262;
end
3082:begin
x_i <= 65416;
end
3083:begin
x_i <= 127;
end
3084:begin
x_i <= 354;
end
3085:begin
x_i <= 289;
end
3086:begin
x_i <= 196;
end
3087:begin
x_i <= 95;
end
3088:begin
x_i <= 65304;
end
3089:begin
x_i <= 65180;
end
3090:begin
x_i <= 65273;
end
3091:begin
x_i <= 65351;
end
3092:begin
x_i <= 65486;
end
3093:begin
x_i <= 204;
end
3094:begin
x_i <= 266;
end
3095:begin
x_i <= 136;
end
3096:begin
x_i <= 81;
end
3097:begin
x_i <= 65456;
end
3098:begin
x_i <= 65243;
end
3099:begin
x_i <= 65224;
end
3100:begin
x_i <= 65302;
end
3101:begin
x_i <= 65415;
end
3102:begin
x_i <= 13;
end
3103:begin
x_i <= 120;
end
3104:begin
x_i <= 87;
end
3105:begin
x_i <= 65507;
end
3106:begin
x_i <= 65406;
end
3107:begin
x_i <= 65295;
end
3108:begin
x_i <= 65246;
end
3109:begin
x_i <= 65394;
end
3110:begin
x_i <= 4;
end
3111:begin
x_i <= 107;
end
3112:begin
x_i <= 164;
end
3113:begin
x_i <= 169;
end
3114:begin
x_i <= 32;
end
3115:begin
x_i <= 65458;
end
3116:begin
x_i <= 65375;
end
3117:begin
x_i <= 65351;
end
3118:begin
x_i <= 65433;
end
3119:begin
x_i <= 24;
end
3120:begin
x_i <= 85;
end
3121:begin
x_i <= 137;
end
3122:begin
x_i <= 210;
end
3123:begin
x_i <= 57;
end
3124:begin
x_i <= 65470;
end
3125:begin
x_i <= 65411;
end
3126:begin
x_i <= 65318;
end
3127:begin
x_i <= 65250;
end
3128:begin
x_i <= 65377;
end
3129:begin
x_i <= 65508;
end
3130:begin
x_i <= 27;
end
3131:begin
x_i <= 43;
end
3132:begin
x_i <= 67;
end
3133:begin
x_i <= 65527;
end
3134:begin
x_i <= 65428;
end
3135:begin
x_i <= 65388;
end
3136:begin
x_i <= 65335;
end
3137:begin
x_i <= 65375;
end
3138:begin
x_i <= 65485;
end
3139:begin
x_i <= 27;
end
3140:begin
x_i <= 87;
end
3141:begin
x_i <= 187;
end
3142:begin
x_i <= 123;
end
3143:begin
x_i <= 3;
end
3144:begin
x_i <= 65485;
end
3145:begin
x_i <= 65458;
end
3146:begin
x_i <= 65374;
end
3147:begin
x_i <= 65410;
end
3148:begin
x_i <= 65534;
end
3149:begin
x_i <= 65524;
end
3150:begin
x_i <= 34;
end
3151:begin
x_i <= 122;
end
3152:begin
x_i <= 66;
end
3153:begin
x_i <= 65509;
end
3154:begin
x_i <= 65451;
end
3155:begin
x_i <= 65472;
end
3156:begin
x_i <= 65421;
end
3157:begin
x_i <= 65467;
end
3158:begin
x_i <= 21;
end
3159:begin
x_i <= 65516;
end
3160:begin
x_i <= 65442;
end
3161:begin
x_i <= 53;
end
3162:begin
x_i <= 65493;
end
3163:begin
x_i <= 65486;
end
3164:begin
x_i <= 32;
end
3165:begin
x_i <= 65532;
end
3166:begin
x_i <= 65532;
end
3167:begin
x_i <= 65454;
end
3168:begin
x_i <= 34;
end
3169:begin
x_i <= 46;
end
3170:begin
x_i <= 12;
end
3171:begin
x_i <= 169;
end
3172:begin
x_i <= 139;
end
3173:begin
x_i <= 66;
end
3174:begin
x_i <= 52;
end
3175:begin
x_i <= 21;
end
3176:begin
x_i <= 65490;
end
3177:begin
x_i <= 65424;
end
3178:begin
x_i <= 65433;
end
3179:begin
x_i <= 65435;
end
3180:begin
x_i <= 65466;
end
3181:begin
x_i <= 65467;
end
3182:begin
x_i <= 65532;
end
3183:begin
x_i <= 37;
end
3184:begin
x_i <= 65520;
end
3185:begin
x_i <= 65480;
end
3186:begin
x_i <= 65458;
end
3187:begin
x_i <= 65484;
end
3188:begin
x_i <= 65471;
end
3189:begin
x_i <= 65457;
end
3190:begin
x_i <= 65534;
end
3191:begin
x_i <= 65522;
end
3192:begin
x_i <= 65479;
end
3193:begin
x_i <= 65519;
end
3194:begin
x_i <= 65502;
end
3195:begin
x_i <= 65487;
end
3196:begin
x_i <= 65475;
end
3197:begin
x_i <= 65532;
end
3198:begin
x_i <= 65515;
end
3199:begin
x_i <= 65508;
end
3200:begin
x_i <= 10;
end
3201:begin
x_i <= 23;
end
3202:begin
x_i <= 65519;
end
3203:begin
x_i <= 65503;
end
3204:begin
x_i <= 65471;
end
3205:begin
x_i <= 65484;
end
3206:begin
x_i <= 65436;
end
3207:begin
x_i <= 65468;
end
3208:begin
x_i <= 65526;
end
3209:begin
x_i <= 1;
end
3210:begin
x_i <= 65524;
end
3211:begin
x_i <= 65505;
end
3212:begin
x_i <= 65506;
end
3213:begin
x_i <= 65496;
end
3214:begin
x_i <= 65450;
end
3215:begin
x_i <= 65507;
end
3216:begin
x_i <= 10;
end
3217:begin
x_i <= 20;
end
3218:begin
x_i <= 65;
end
3219:begin
x_i <= 120;
end
3220:begin
x_i <= 140;
end
3221:begin
x_i <= 58;
end
3222:begin
x_i <= 65519;
end
3223:begin
x_i <= 65513;
end
3224:begin
x_i <= 65444;
end
3225:begin
x_i <= 65470;
end
3226:begin
x_i <= 65512;
end
3227:begin
x_i <= 40;
end
3228:begin
x_i <= 67;
end
3229:begin
x_i <= 66;
end
3230:begin
x_i <= 52;
end
3231:begin
x_i <= 1;
end
3232:begin
x_i <= 65491;
end
3233:begin
x_i <= 65471;
end
3234:begin
x_i <= 65458;
end
3235:begin
x_i <= 65509;
end
3236:begin
x_i <= 65499;
end
3237:begin
x_i <= 65474;
end
3238:begin
x_i <= 29;
end
3239:begin
x_i <= 65534;
end
3240:begin
x_i <= 65497;
end
3241:begin
x_i <= 65532;
end
3242:begin
x_i <= 65519;
end
3243:begin
x_i <= 65464;
end
3244:begin
x_i <= 65468;
end
3245:begin
x_i <= 65510;
end
3246:begin
x_i <= 65509;
end
3247:begin
x_i <= 65476;
end
3248:begin
x_i <= 65506;
end
3249:begin
x_i <= 65508;
end
3250:begin
x_i <= 17;
end
3251:begin
x_i <= 18;
end
3252:begin
x_i <= 22;
end
3253:begin
x_i <= 3;
end
3254:begin
x_i <= 65492;
end
3255:begin
x_i <= 65495;
end
3256:begin
x_i <= 65488;
end
3257:begin
x_i <= 65477;
end
3258:begin
x_i <= 16;
end
3259:begin
x_i <= 65524;
end
3260:begin
x_i <= 44;
end
3261:begin
x_i <= 80;
end
3262:begin
x_i <= 29;
end
3263:begin
x_i <= 65514;
end
3264:begin
x_i <= 65407;
end
3265:begin
x_i <= 65441;
end
3266:begin
x_i <= 65423;
end
3267:begin
x_i <= 65443;
end
3268:begin
x_i <= 17;
end
3269:begin
x_i <= 35;
end
3270:begin
x_i <= 64;
end
3271:begin
x_i <= 54;
end
3272:begin
x_i <= 33;
end
3273:begin
x_i <= 65478;
end
3274:begin
x_i <= 65471;
end
3275:begin
x_i <= 65488;
end
3276:begin
x_i <= 65476;
end
3277:begin
x_i <= 65487;
end
3278:begin
x_i <= 0;
end
3279:begin
x_i <= 65481;
end
3280:begin
x_i <= 65483;
end
3281:begin
x_i <= 65476;
end
3282:begin
x_i <= 65495;
end
3283:begin
x_i <= 65495;
end
3284:begin
x_i <= 65517;
end
3285:begin
x_i <= 8;
end
3286:begin
x_i <= 65513;
end
3287:begin
x_i <= 65435;
end
3288:begin
x_i <= 65500;
end
3289:begin
x_i <= 0;
end
3290:begin
x_i <= 65526;
end
3291:begin
x_i <= 31;
end
3292:begin
x_i <= 65533;
end
3293:begin
x_i <= 65475;
end
3294:begin
x_i <= 65470;
end
3295:begin
x_i <= 65432;
end
3296:begin
x_i <= 65434;
end
3297:begin
x_i <= 65446;
end
3298:begin
x_i <= 65473;
end
3299:begin
x_i <= 65514;
end
3300:begin
x_i <= 65530;
end
3301:begin
x_i <= 65499;
end
3302:begin
x_i <= 74;
end
3303:begin
x_i <= 59;
end
3304:begin
x_i <= 65483;
end
3305:begin
x_i <= 65535;
end
3306:begin
x_i <= 65524;
end
3307:begin
x_i <= 65457;
end
3308:begin
x_i <= 65507;
end
3309:begin
x_i <= 17;
end
3310:begin
x_i <= 47;
end
3311:begin
x_i <= 7;
end
3312:begin
x_i <= 2;
end
3313:begin
x_i <= 59;
end
3314:begin
x_i <= 65528;
end
3315:begin
x_i <= 65481;
end
3316:begin
x_i <= 65497;
end
3317:begin
x_i <= 65468;
end
3318:begin
x_i <= 65438;
end
3319:begin
x_i <= 65507;
end
3320:begin
x_i <= 3;
end
3321:begin
x_i <= 65530;
end
3322:begin
x_i <= 94;
end
3323:begin
x_i <= 93;
end
3324:begin
x_i <= 16;
end
3325:begin
x_i <= 65503;
end
3326:begin
x_i <= 65477;
end
3327:begin
x_i <= 65426;
end
3328:begin
x_i <= 65424;
end
3329:begin
x_i <= 65486;
end
3330:begin
x_i <= 65533;
end
3331:begin
x_i <= 65517;
end
3332:begin
x_i <= 25;
end
3333:begin
x_i <= 30;
end
3334:begin
x_i <= 65510;
end
3335:begin
x_i <= 65483;
end
3336:begin
x_i <= 65479;
end
3337:begin
x_i <= 65445;
end
3338:begin
x_i <= 65403;
end
3339:begin
x_i <= 65490;
end
3340:begin
x_i <= 23;
end
3341:begin
x_i <= 0;
end
3342:begin
x_i <= 65535;
end
3343:begin
x_i <= 65531;
end
3344:begin
x_i <= 65535;
end
3345:begin
x_i <= 65443;
end
3346:begin
x_i <= 65464;
end
3347:begin
x_i <= 8;
end
3348:begin
x_i <= 65520;
end
3349:begin
x_i <= 16;
end
3350:begin
x_i <= 110;
end
3351:begin
x_i <= 100;
end
3352:begin
x_i <= 65528;
end
3353:begin
x_i <= 65488;
end
3354:begin
x_i <= 65485;
end
3355:begin
x_i <= 65488;
end
3356:begin
x_i <= 65446;
end
3357:begin
x_i <= 13;
end
3358:begin
x_i <= 45;
end
3359:begin
x_i <= 11;
end
3360:begin
x_i <= 44;
end
3361:begin
x_i <= 104;
end
3362:begin
x_i <= 65516;
end
3363:begin
x_i <= 65484;
end
3364:begin
x_i <= 65475;
end
3365:begin
x_i <= 65446;
end
3366:begin
x_i <= 65420;
end
3367:begin
x_i <= 65494;
end
3368:begin
x_i <= 60;
end
3369:begin
x_i <= 32;
end
3370:begin
x_i <= 8;
end
3371:begin
x_i <= 56;
end
3372:begin
x_i <= 65471;
end
3373:begin
x_i <= 65465;
end
3374:begin
x_i <= 65481;
end
3375:begin
x_i <= 65466;
end
3376:begin
x_i <= 65481;
end
3377:begin
x_i <= 3;
end
3378:begin
x_i <= 45;
end
3379:begin
x_i <= 65523;
end
3380:begin
x_i <= 17;
end
3381:begin
x_i <= 17;
end
3382:begin
x_i <= 65449;
end
3383:begin
x_i <= 65499;
end
3384:begin
x_i <= 65462;
end
3385:begin
x_i <= 65520;
end
3386:begin
x_i <= 65481;
end
3387:begin
x_i <= 38;
end
3388:begin
x_i <= 34;
end
3389:begin
x_i <= 65496;
end
3390:begin
x_i <= 65505;
end
3391:begin
x_i <= 65483;
end
3392:begin
x_i <= 65485;
end
3393:begin
x_i <= 65497;
end
3394:begin
x_i <= 15;
end
3395:begin
x_i <= 62;
end
3396:begin
x_i <= 49;
end
3397:begin
x_i <= 86;
end
3398:begin
x_i <= 56;
end
3399:begin
x_i <= 65512;
end
3400:begin
x_i <= 65469;
end
3401:begin
x_i <= 65427;
end
3402:begin
x_i <= 65450;
end
3403:begin
x_i <= 1;
end
3404:begin
x_i <= 32;
end
3405:begin
x_i <= 113;
end
3406:begin
x_i <= 16;
end
3407:begin
x_i <= 23;
end
3408:begin
x_i <= 14;
end
3409:begin
x_i <= 65450;
end
3410:begin
x_i <= 65491;
end
3411:begin
x_i <= 65523;
end
3412:begin
x_i <= 65494;
end
3413:begin
x_i <= 69;
end
3414:begin
x_i <= 37;
end
3415:begin
x_i <= 40;
end
3416:begin
x_i <= 109;
end
3417:begin
x_i <= 77;
end
3418:begin
x_i <= 24;
end
3419:begin
x_i <= 65516;
end
3420:begin
x_i <= 65486;
end
3421:begin
x_i <= 65446;
end
3422:begin
x_i <= 65463;
end
3423:begin
x_i <= 65520;
end
3424:begin
x_i <= 19;
end
3425:begin
x_i <= 65499;
end
3426:begin
x_i <= 65520;
end
3427:begin
x_i <= 65523;
end
3428:begin
x_i <= 65520;
end
3429:begin
x_i <= 34;
end
3430:begin
x_i <= 66;
end
3431:begin
x_i <= 49;
end
3432:begin
x_i <= 65533;
end
3433:begin
x_i <= 34;
end
3434:begin
x_i <= 25;
end
3435:begin
x_i <= 65499;
end
3436:begin
x_i <= 8;
end
3437:begin
x_i <= 65510;
end
3438:begin
x_i <= 65523;
end
3439:begin
x_i <= 1;
end
3440:begin
x_i <= 6;
end
3441:begin
x_i <= 40;
end
3442:begin
x_i <= 65520;
end
3443:begin
x_i <= 65507;
end
3444:begin
x_i <= 33;
end
3445:begin
x_i <= 23;
end
3446:begin
x_i <= 0;
end
3447:begin
x_i <= 1;
end
3448:begin
x_i <= 65468;
end
3449:begin
x_i <= 65464;
end
3450:begin
x_i <= 65503;
end
3451:begin
x_i <= 2;
end
3452:begin
x_i <= 1;
end
3453:begin
x_i <= 65465;
end
3454:begin
x_i <= 65418;
end
3455:begin
x_i <= 65389;
end
3456:begin
x_i <= 65473;
end
3457:begin
x_i <= 17;
end
3458:begin
x_i <= 65513;
end
3459:begin
x_i <= 65508;
end
3460:begin
x_i <= 65435;
end
3461:begin
x_i <= 65454;
end
3462:begin
x_i <= 65501;
end
3463:begin
x_i <= 65415;
end
3464:begin
x_i <= 65497;
end
3465:begin
x_i <= 65450;
end
3466:begin
x_i <= 65427;
end
3467:begin
x_i <= 65419;
end
3468:begin
x_i <= 65380;
end
3469:begin
x_i <= 65434;
end
3470:begin
x_i <= 65395;
end
3471:begin
x_i <= 65393;
end
3472:begin
x_i <= 65432;
end
3473:begin
x_i <= 65501;
end
3474:begin
x_i <= 65470;
end
3475:begin
x_i <= 65472;
end
3476:begin
x_i <= 65475;
end
3477:begin
x_i <= 65420;
end
3478:begin
x_i <= 65440;
end
3479:begin
x_i <= 65425;
end
3480:begin
x_i <= 65450;
end
3481:begin
x_i <= 65424;
end
3482:begin
x_i <= 65387;
end
3483:begin
x_i <= 65460;
end
3484:begin
x_i <= 65467;
end
3485:begin
x_i <= 65522;
end
3486:begin
x_i <= 65516;
end
3487:begin
x_i <= 65534;
end
3488:begin
x_i <= 65524;
end
3489:begin
x_i <= 65500;
end
3490:begin
x_i <= 65512;
end
3491:begin
x_i <= 28;
end
3492:begin
x_i <= 21;
end
3493:begin
x_i <= 38;
end
3494:begin
x_i <= 100;
end
3495:begin
x_i <= 106;
end
3496:begin
x_i <= 55;
end
3497:begin
x_i <= 25;
end
3498:begin
x_i <= 35;
end
3499:begin
x_i <= 65522;
end
3500:begin
x_i <= 43;
end
3501:begin
x_i <= 40;
end
3502:begin
x_i <= 104;
end
3503:begin
x_i <= 122;
end
3504:begin
x_i <= 94;
end
3505:begin
x_i <= 151;
end
3506:begin
x_i <= 88;
end
3507:begin
x_i <= 111;
end
3508:begin
x_i <= 113;
end
3509:begin
x_i <= 54;
end
3510:begin
x_i <= 122;
end
3511:begin
x_i <= 116;
end
3512:begin
x_i <= 190;
end
3513:begin
x_i <= 250;
end
3514:begin
x_i <= 269;
end
3515:begin
x_i <= 232;
end
3516:begin
x_i <= 193;
end
3517:begin
x_i <= 136;
end
3518:begin
x_i <= 81;
end
3519:begin
x_i <= 92;
end
3520:begin
x_i <= 89;
end
3521:begin
x_i <= 176;
end
3522:begin
x_i <= 124;
end
3523:begin
x_i <= 175;
end
3524:begin
x_i <= 275;
end
3525:begin
x_i <= 326;
end
3526:begin
x_i <= 238;
end
3527:begin
x_i <= 161;
end
3528:begin
x_i <= 52;
end
3529:begin
x_i <= 65446;
end
3530:begin
x_i <= 65298;
end
3531:begin
x_i <= 65327;
end
3532:begin
x_i <= 65384;
end
3533:begin
x_i <= 65369;
end
3534:begin
x_i <= 65412;
end
3535:begin
x_i <= 65495;
end
3536:begin
x_i <= 2;
end
3537:begin
x_i <= 65367;
end
3538:begin
x_i <= 65344;
end
3539:begin
x_i <= 65365;
end
3540:begin
x_i <= 65172;
end
3541:begin
x_i <= 65108;
end
3542:begin
x_i <= 65243;
end
3543:begin
x_i <= 65328;
end
3544:begin
x_i <= 65379;
end
3545:begin
x_i <= 65490;
end
3546:begin
x_i <= 65525;
end
3547:begin
x_i <= 65518;
end
3548:begin
x_i <= 65339;
end
3549:begin
x_i <= 65249;
end
3550:begin
x_i <= 65203;
end
3551:begin
x_i <= 65138;
end
3552:begin
x_i <= 65174;
end
3553:begin
x_i <= 65249;
end
3554:begin
x_i <= 65323;
end
3555:begin
x_i <= 65413;
end
3556:begin
x_i <= 65459;
end
3557:begin
x_i <= 65440;
end
3558:begin
x_i <= 65418;
end
3559:begin
x_i <= 65321;
end
3560:begin
x_i <= 65209;
end
3561:begin
x_i <= 65177;
end
3562:begin
x_i <= 65211;
end
3563:begin
x_i <= 65243;
end
3564:begin
x_i <= 65331;
end
3565:begin
x_i <= 65395;
end
3566:begin
x_i <= 65479;
end
3567:begin
x_i <= 65471;
end
3568:begin
x_i <= 65466;
end
3569:begin
x_i <= 65495;
end
3570:begin
x_i <= 65428;
end
3571:begin
x_i <= 65422;
end
3572:begin
x_i <= 65433;
end
3573:begin
x_i <= 65505;
end
3574:begin
x_i <= 65525;
end
3575:begin
x_i <= 4;
end
3576:begin
x_i <= 25;
end
3577:begin
x_i <= 55;
end
3578:begin
x_i <= 65530;
end
3579:begin
x_i <= 65493;
end
3580:begin
x_i <= 65526;
end
3581:begin
x_i <= 65525;
end
3582:begin
x_i <= 65521;
end
3583:begin
x_i <= 32;
end
3584:begin
x_i <= 95;
end
3585:begin
x_i <= 125;
end
3586:begin
x_i <= 79;
end
3587:begin
x_i <= 91;
end
3588:begin
x_i <= 90;
end
3589:begin
x_i <= 72;
end
3590:begin
x_i <= 65534;
end
3591:begin
x_i <= 4;
end
3592:begin
x_i <= 82;
end
3593:begin
x_i <= 138;
end
3594:begin
x_i <= 234;
end
3595:begin
x_i <= 338;
end
3596:begin
x_i <= 401;
end
3597:begin
x_i <= 264;
end
3598:begin
x_i <= 206;
end
3599:begin
x_i <= 139;
end
3600:begin
x_i <= 54;
end
3601:begin
x_i <= 52;
end
3602:begin
x_i <= 65527;
end
3603:begin
x_i <= 155;
end
3604:begin
x_i <= 252;
end
3605:begin
x_i <= 270;
end
3606:begin
x_i <= 362;
end
3607:begin
x_i <= 441;
end
3608:begin
x_i <= 288;
end
3609:begin
x_i <= 78;
end
3610:begin
x_i <= 65505;
end
3611:begin
x_i <= 65437;
end
3612:begin
x_i <= 65262;
end
3613:begin
x_i <= 65207;
end
3614:begin
x_i <= 65314;
end
3615:begin
x_i <= 65438;
end
3616:begin
x_i <= 65395;
end
3617:begin
x_i <= 34;
end
3618:begin
x_i <= 141;
end
3619:begin
x_i <= 39;
end
3620:begin
x_i <= 65452;
end
3621:begin
x_i <= 65295;
end
3622:begin
x_i <= 65250;
end
3623:begin
x_i <= 65270;
end
3624:begin
x_i <= 65290;
end
3625:begin
x_i <= 65485;
end
3626:begin
x_i <= 65534;
end
3627:begin
x_i <= 52;
end
3628:begin
x_i <= 5;
end
3629:begin
x_i <= 65506;
end
3630:begin
x_i <= 65522;
end
3631:begin
x_i <= 65383;
end
3632:begin
x_i <= 65190;
end
3633:begin
x_i <= 65128;
end
3634:begin
x_i <= 65165;
end
3635:begin
x_i <= 65198;
end
3636:begin
x_i <= 65321;
end
3637:begin
x_i <= 65424;
end
3638:begin
x_i <= 65496;
end
3639:begin
x_i <= 65466;
end
3640:begin
x_i <= 65387;
end
3641:begin
x_i <= 65436;
end
3642:begin
x_i <= 65327;
end
3643:begin
x_i <= 65233;
end
3644:begin
x_i <= 65275;
end
3645:begin
x_i <= 65264;
end
3646:begin
x_i <= 65335;
end
3647:begin
x_i <= 65397;
end
3648:begin
x_i <= 65424;
end
3649:begin
x_i <= 65472;
end
3650:begin
x_i <= 65453;
end
3651:begin
x_i <= 65397;
end
3652:begin
x_i <= 65466;
end
3653:begin
x_i <= 65490;
end
3654:begin
x_i <= 2;
end
3655:begin
x_i <= 10;
end
3656:begin
x_i <= 13;
end
3657:begin
x_i <= 55;
end
3658:begin
x_i <= 65516;
end
3659:begin
x_i <= 65507;
end
3660:begin
x_i <= 65466;
end
3661:begin
x_i <= 65397;
end
3662:begin
x_i <= 65403;
end
3663:begin
x_i <= 65427;
end
3664:begin
x_i <= 65500;
end
3665:begin
x_i <= 65532;
end
3666:begin
x_i <= 35;
end
3667:begin
x_i <= 47;
end
3668:begin
x_i <= 101;
end
3669:begin
x_i <= 135;
end
3670:begin
x_i <= 135;
end
3671:begin
x_i <= 133;
end
3672:begin
x_i <= 47;
end
3673:begin
x_i <= 65506;
end
3674:begin
x_i <= 65529;
end
3675:begin
x_i <= 49;
end
3676:begin
x_i <= 88;
end
3677:begin
x_i <= 109;
end
3678:begin
x_i <= 209;
end
3679:begin
x_i <= 173;
end
3680:begin
x_i <= 123;
end
3681:begin
x_i <= 172;
end
3682:begin
x_i <= 119;
end
3683:begin
x_i <= 166;
end
3684:begin
x_i <= 127;
end
3685:begin
x_i <= 240;
end
3686:begin
x_i <= 371;
end
3687:begin
x_i <= 394;
end
3688:begin
x_i <= 440;
end
3689:begin
x_i <= 399;
end
3690:begin
x_i <= 318;
end
3691:begin
x_i <= 215;
end
3692:begin
x_i <= 29;
end
3693:begin
x_i <= 15;
end
3694:begin
x_i <= 1;
end
3695:begin
x_i <= 65436;
end
3696:begin
x_i <= 65396;
end
3697:begin
x_i <= 65493;
end
3698:begin
x_i <= 65489;
end
3699:begin
x_i <= 65421;
end
3700:begin
x_i <= 65423;
end
3701:begin
x_i <= 65445;
end
3702:begin
x_i <= 65442;
end
3703:begin
x_i <= 65322;
end
3704:begin
x_i <= 65419;
end
3705:begin
x_i <= 65513;
end
3706:begin
x_i <= 65449;
end
3707:begin
x_i <= 65431;
end
3708:begin
x_i <= 65493;
end
3709:begin
x_i <= 65445;
end
3710:begin
x_i <= 65428;
end
3711:begin
x_i <= 65422;
end
3712:begin
x_i <= 65453;
end
3713:begin
x_i <= 65432;
end
3714:begin
x_i <= 65337;
end
3715:begin
x_i <= 65368;
end
3716:begin
x_i <= 65395;
end
3717:begin
x_i <= 65417;
end
3718:begin
x_i <= 65422;
end
3719:begin
x_i <= 65443;
end
3720:begin
x_i <= 65480;
end
3721:begin
x_i <= 65446;
end
3722:begin
x_i <= 65362;
end
3723:begin
x_i <= 65301;
end
3724:begin
x_i <= 65312;
end
3725:begin
x_i <= 65244;
end
3726:begin
x_i <= 65223;
end
3727:begin
x_i <= 65274;
end
3728:begin
x_i <= 65283;
end
3729:begin
x_i <= 65299;
end
3730:begin
x_i <= 65379;
end
3731:begin
x_i <= 65447;
end
3732:begin
x_i <= 65422;
end
3733:begin
x_i <= 65397;
end
3734:begin
x_i <= 65442;
end
3735:begin
x_i <= 65490;
end
3736:begin
x_i <= 65484;
end
3737:begin
x_i <= 65460;
end
3738:begin
x_i <= 5;
end
3739:begin
x_i <= 0;
end
3740:begin
x_i <= 65504;
end
3741:begin
x_i <= 65480;
end
3742:begin
x_i <= 65491;
end
3743:begin
x_i <= 65478;
end
3744:begin
x_i <= 65444;
end
3745:begin
x_i <= 65464;
end
3746:begin
x_i <= 65512;
end
3747:begin
x_i <= 65493;
end
3748:begin
x_i <= 65505;
end
3749:begin
x_i <= 65478;
end
3750:begin
x_i <= 65488;
end
3751:begin
x_i <= 65479;
end
3752:begin
x_i <= 65455;
end
3753:begin
x_i <= 65475;
end
3754:begin
x_i <= 65510;
end
3755:begin
x_i <= 36;
end
3756:begin
x_i <= 53;
end
3757:begin
x_i <= 99;
end
3758:begin
x_i <= 63;
end
3759:begin
x_i <= 56;
end
3760:begin
x_i <= 86;
end
3761:begin
x_i <= 79;
end
3762:begin
x_i <= 36;
end
3763:begin
x_i <= 20;
end
3764:begin
x_i <= 77;
end
3765:begin
x_i <= 110;
end
3766:begin
x_i <= 130;
end
3767:begin
x_i <= 117;
end
3768:begin
x_i <= 160;
end
3769:begin
x_i <= 230;
end
3770:begin
x_i <= 177;
end
3771:begin
x_i <= 133;
end
3772:begin
x_i <= 138;
end
3773:begin
x_i <= 112;
end
3774:begin
x_i <= 115;
end
3775:begin
x_i <= 28;
end
3776:begin
x_i <= 141;
end
3777:begin
x_i <= 152;
end
3778:begin
x_i <= 145;
end
3779:begin
x_i <= 279;
end
3780:begin
x_i <= 346;
end
3781:begin
x_i <= 389;
end
3782:begin
x_i <= 288;
end
3783:begin
x_i <= 129;
end
3784:begin
x_i <= 59;
end
3785:begin
x_i <= 65492;
end
3786:begin
x_i <= 65417;
end
3787:begin
x_i <= 65364;
end
3788:begin
x_i <= 65425;
end
3789:begin
x_i <= 65431;
end
3790:begin
x_i <= 65438;
end
3791:begin
x_i <= 65504;
end
3792:begin
x_i <= 41;
end
3793:begin
x_i <= 71;
end
3794:begin
x_i <= 10;
end
3795:begin
x_i <= 65462;
end
3796:begin
x_i <= 65416;
end
3797:begin
x_i <= 65323;
end
3798:begin
x_i <= 65335;
end
3799:begin
x_i <= 65372;
end
3800:begin
x_i <= 65456;
end
3801:begin
x_i <= 1;
end
3802:begin
x_i <= 38;
end
3803:begin
x_i <= 50;
end
3804:begin
x_i <= 65535;
end
3805:begin
x_i <= 65461;
end
3806:begin
x_i <= 65378;
end
3807:begin
x_i <= 65304;
end
3808:begin
x_i <= 65275;
end
3809:begin
x_i <= 65278;
end
3810:begin
x_i <= 65321;
end
3811:begin
x_i <= 65418;
end
3812:begin
x_i <= 65455;
end
3813:begin
x_i <= 65493;
end
3814:begin
x_i <= 65506;
end
3815:begin
x_i <= 65493;
end
3816:begin
x_i <= 65414;
end
3817:begin
x_i <= 65297;
end
3818:begin
x_i <= 65220;
end
3819:begin
x_i <= 65202;
end
3820:begin
x_i <= 65178;
end
3821:begin
x_i <= 65279;
end
3822:begin
x_i <= 65376;
end
3823:begin
x_i <= 65491;
end
3824:begin
x_i <= 65517;
end
3825:begin
x_i <= 22;
end
3826:begin
x_i <= 22;
end
3827:begin
x_i <= 65493;
end
3828:begin
x_i <= 65442;
end
3829:begin
x_i <= 65455;
end
3830:begin
x_i <= 65442;
end
3831:begin
x_i <= 65428;
end
3832:begin
x_i <= 65419;
end
3833:begin
x_i <= 65462;
end
3834:begin
x_i <= 65494;
end
3835:begin
x_i <= 65485;
end
3836:begin
x_i <= 65495;
end
3837:begin
x_i <= 65515;
end
3838:begin
x_i <= 65508;
end
3839:begin
x_i <= 65492;
end
3840:begin
x_i <= 65452;
end
3841:begin
x_i <= 65472;
end
3842:begin
x_i <= 65473;
end
3843:begin
x_i <= 65494;
end
3844:begin
x_i <= 65528;
end
3845:begin
x_i <= 39;
end
3846:begin
x_i <= 83;
end
3847:begin
x_i <= 112;
end
3848:begin
x_i <= 104;
end
3849:begin
x_i <= 122;
end
3850:begin
x_i <= 97;
end
3851:begin
x_i <= 80;
end
3852:begin
x_i <= 28;
end
3853:begin
x_i <= 7;
end
3854:begin
x_i <= 65524;
end
3855:begin
x_i <= 65527;
end
3856:begin
x_i <= 3;
end
3857:begin
x_i <= 109;
end
3858:begin
x_i <= 202;
end
3859:begin
x_i <= 264;
end
3860:begin
x_i <= 249;
end
3861:begin
x_i <= 239;
end
3862:begin
x_i <= 195;
end
3863:begin
x_i <= 190;
end
3864:begin
x_i <= 151;
end
3865:begin
x_i <= 66;
end
3866:begin
x_i <= 52;
end
3867:begin
x_i <= 95;
end
3868:begin
x_i <= 45;
end
3869:begin
x_i <= 88;
end
3870:begin
x_i <= 188;
end
3871:begin
x_i <= 237;
end
3872:begin
x_i <= 250;
end
3873:begin
x_i <= 168;
end
3874:begin
x_i <= 35;
end
3875:begin
x_i <= 65525;
end
3876:begin
x_i <= 65461;
end
3877:begin
x_i <= 65482;
end
3878:begin
x_i <= 65484;
end
3879:begin
x_i <= 65459;
end
3880:begin
x_i <= 65472;
end
3881:begin
x_i <= 65397;
end
3882:begin
x_i <= 65400;
end
3883:begin
x_i <= 65424;
end
3884:begin
x_i <= 65410;
end
3885:begin
x_i <= 65404;
end
3886:begin
x_i <= 65445;
end
3887:begin
x_i <= 65495;
end
3888:begin
x_i <= 65486;
end
3889:begin
x_i <= 65487;
end
3890:begin
x_i <= 8;
end
3891:begin
x_i <= 8;
end
3892:begin
x_i <= 65505;
end
3893:begin
x_i <= 65463;
end
3894:begin
x_i <= 65475;
end
3895:begin
x_i <= 65497;
end
3896:begin
x_i <= 65466;
end
3897:begin
x_i <= 65402;
end
3898:begin
x_i <= 65377;
end
3899:begin
x_i <= 65414;
end
3900:begin
x_i <= 65402;
end
3901:begin
x_i <= 65458;
end
3902:begin
x_i <= 65460;
end
3903:begin
x_i <= 65403;
end
3904:begin
x_i <= 65343;
end
3905:begin
x_i <= 65340;
end
3906:begin
x_i <= 65398;
end
3907:begin
x_i <= 65410;
end
3908:begin
x_i <= 65428;
end
3909:begin
x_i <= 65436;
end
3910:begin
x_i <= 65456;
end
3911:begin
x_i <= 65423;
end
3912:begin
x_i <= 65420;
end
3913:begin
x_i <= 65416;
end
3914:begin
x_i <= 65399;
end
3915:begin
x_i <= 65378;
end
3916:begin
x_i <= 65406;
end
3917:begin
x_i <= 65458;
end
3918:begin
x_i <= 65506;
end
3919:begin
x_i <= 65531;
end
3920:begin
x_i <= 31;
end
3921:begin
x_i <= 25;
end
3922:begin
x_i <= 21;
end
3923:begin
x_i <= 65503;
end
3924:begin
x_i <= 65489;
end
3925:begin
x_i <= 65441;
end
3926:begin
x_i <= 65409;
end
3927:begin
x_i <= 65420;
end
3928:begin
x_i <= 65449;
end
3929:begin
x_i <= 65499;
end
3930:begin
x_i <= 65527;
end
3931:begin
x_i <= 65526;
end
3932:begin
x_i <= 2;
end
3933:begin
x_i <= 65521;
end
3934:begin
x_i <= 65487;
end
3935:begin
x_i <= 65508;
end
3936:begin
x_i <= 65507;
end
3937:begin
x_i <= 9;
end
3938:begin
x_i <= 31;
end
3939:begin
x_i <= 30;
end
3940:begin
x_i <= 103;
end
3941:begin
x_i <= 79;
end
3942:begin
x_i <= 38;
end
3943:begin
x_i <= 13;
end
3944:begin
x_i <= 36;
end
3945:begin
x_i <= 33;
end
3946:begin
x_i <= 18;
end
3947:begin
x_i <= 7;
end
3948:begin
x_i <= 90;
end
3949:begin
x_i <= 79;
end
3950:begin
x_i <= 21;
end
3951:begin
x_i <= 37;
end
3952:begin
x_i <= 53;
end
3953:begin
x_i <= 103;
end
3954:begin
x_i <= 88;
end
3955:begin
x_i <= 152;
end
3956:begin
x_i <= 212;
end
3957:begin
x_i <= 183;
end
3958:begin
x_i <= 197;
end
3959:begin
x_i <= 145;
end
3960:begin
x_i <= 122;
end
3961:begin
x_i <= 91;
end
3962:begin
x_i <= 65532;
end
3963:begin
x_i <= 43;
end
3964:begin
x_i <= 88;
end
3965:begin
x_i <= 88;
end
3966:begin
x_i <= 197;
end
3967:begin
x_i <= 223;
end
3968:begin
x_i <= 249;
end
3969:begin
x_i <= 177;
end
3970:begin
x_i <= 118;
end
3971:begin
x_i <= 30;
end
3972:begin
x_i <= 65357;
end
3973:begin
x_i <= 65220;
end
3974:begin
x_i <= 65267;
end
3975:begin
x_i <= 65256;
end
3976:begin
x_i <= 65291;
end
3977:begin
x_i <= 65413;
end
3978:begin
x_i <= 46;
end
3979:begin
x_i <= 73;
end
3980:begin
x_i <= 65;
end
3981:begin
x_i <= 89;
end
3982:begin
x_i <= 21;
end
3983:begin
x_i <= 65448;
end
3984:begin
x_i <= 65350;
end
3985:begin
x_i <= 65387;
end
3986:begin
x_i <= 65443;
end
3987:begin
x_i <= 65462;
end
3988:begin
x_i <= 27;
end
3989:begin
x_i <= 77;
end
3990:begin
x_i <= 84;
end
3991:begin
x_i <= 37;
end
3992:begin
x_i <= 65466;
end
3993:begin
x_i <= 65443;
end
3994:begin
x_i <= 65381;
end
3995:begin
x_i <= 65351;
end
3996:begin
x_i <= 65396;
end
3997:begin
x_i <= 65454;
end
3998:begin
x_i <= 65489;
end
3999:begin
x_i <= 16;
end
4000:begin
x_i <= 75;
end
4001:begin
x_i <= 37;
end
4002:begin
x_i <= 65484;
end
4003:begin
x_i <= 65373;
end
4004:begin
x_i <= 65315;
end
4005:begin
x_i <= 65286;
end
4006:begin
x_i <= 65319;
end
4007:begin
x_i <= 65358;
end
4008:begin
x_i <= 65429;
end
4009:begin
x_i <= 65493;
end
4010:begin
x_i <= 65504;
end
4011:begin
x_i <= 65491;
end
4012:begin
x_i <= 65495;
end
4013:begin
x_i <= 65494;
end
4014:begin
x_i <= 65450;
end
4015:begin
x_i <= 65452;
end
4016:begin
x_i <= 65412;
end
4017:begin
x_i <= 65396;
end
4018:begin
x_i <= 65368;
end
4019:begin
x_i <= 65417;
end
4020:begin
x_i <= 65393;
end
4021:begin
x_i <= 65379;
end
4022:begin
x_i <= 65401;
end
4023:begin
x_i <= 65406;
end
4024:begin
x_i <= 65400;
end
4025:begin
x_i <= 65432;
end
4026:begin
x_i <= 65429;
end
4027:begin
x_i <= 65441;
end
4028:begin
x_i <= 65526;
end
4029:begin
x_i <= 65525;
end
4030:begin
x_i <= 30;
end
4031:begin
x_i <= 12;
end
4032:begin
x_i <= 65529;
end
4033:begin
x_i <= 65506;
end
4034:begin
x_i <= 65472;
end
4035:begin
x_i <= 65479;
end
4036:begin
x_i <= 65484;
end
4037:begin
x_i <= 65497;
end
4038:begin
x_i <= 7;
end
4039:begin
x_i <= 36;
end
4040:begin
x_i <= 37;
end
4041:begin
x_i <= 32;
end
4042:begin
x_i <= 41;
end
4043:begin
x_i <= 29;
end
4044:begin
x_i <= 6;
end
4045:begin
x_i <= 65531;
end
4046:begin
x_i <= 42;
end
4047:begin
x_i <= 20;
end
4048:begin
x_i <= 34;
end
4049:begin
x_i <= 60;
end
4050:begin
x_i <= 44;
end
4051:begin
x_i <= 40;
end
4052:begin
x_i <= 69;
end
4053:begin
x_i <= 57;
end
4054:begin
x_i <= 104;
end
4055:begin
x_i <= 107;
end
4056:begin
x_i <= 148;
end
4057:begin
x_i <= 250;
end
4058:begin
x_i <= 242;
end
4059:begin
x_i <= 266;
end
4060:begin
x_i <= 250;
end
4061:begin
x_i <= 222;
end
4062:begin
x_i <= 195;
end
4063:begin
x_i <= 199;
end
4064:begin
x_i <= 239;
end
4065:begin
x_i <= 269;
end
4066:begin
x_i <= 158;
end
4067:begin
x_i <= 69;
end
4068:begin
x_i <= 65514;
end
4069:begin
x_i <= 65461;
end
4070:begin
x_i <= 65403;
end
4071:begin
x_i <= 65366;
end
4072:begin
x_i <= 65368;
end
4073:begin
x_i <= 65404;
end
4074:begin
x_i <= 65394;
end
4075:begin
x_i <= 65508;
end
4076:begin
x_i <= 82;
end
4077:begin
x_i <= 30;
end
4078:begin
x_i <= 13;
end
4079:begin
x_i <= 65499;
end
4080:begin
x_i <= 65477;
end
4081:begin
x_i <= 65431;
end
4082:begin
x_i <= 65457;
end
4083:begin
x_i <= 65470;
end
4084:begin
x_i <= 65467;
end
4085:begin
x_i <= 65484;
end
4086:begin
x_i <= 11;
end
4087:begin
x_i <= 10;
end
4088:begin
x_i <= 22;
end
4089:begin
x_i <= 65532;
end
4090:begin
x_i <= 65482;
end
4091:begin
x_i <= 65470;
end
4092:begin
x_i <= 65467;
end
4093:begin
x_i <= 65466;
end
4094:begin
x_i <= 65483;
end
4095:begin
x_i <= 65463;
end
4096:begin
x_i <= 65468;
end
4097:begin
x_i <= 65467;
end
4098:begin
x_i <= 65487;
end
4099:begin
x_i <= 65487;
end
4100:begin
x_i <= 65432;
end
4101:begin
x_i <= 65331;
end
4102:begin
x_i <= 65335;
end
4103:begin
x_i <= 65352;
end
4104:begin
x_i <= 65396;
end
4105:begin
x_i <= 65406;
end
4106:begin
x_i <= 65432;
end
4107:begin
x_i <= 65492;
end
4108:begin
x_i <= 65522;
end
4109:begin
x_i <= 20;
end
4110:begin
x_i <= 32;
end
4111:begin
x_i <= 65507;
end
4112:begin
x_i <= 65431;
end
4113:begin
x_i <= 65416;
end
4114:begin
x_i <= 65375;
end
4115:begin
x_i <= 65337;
end
4116:begin
x_i <= 65348;
end
4117:begin
x_i <= 65320;
end
4118:begin
x_i <= 65344;
end
4119:begin
x_i <= 65383;
end
4120:begin
x_i <= 65455;
end
4121:begin
x_i <= 65430;
end
4122:begin
x_i <= 65446;
end
4123:begin
x_i <= 65440;
end
4124:begin
x_i <= 65393;
end
4125:begin
x_i <= 65363;
end
4126:begin
x_i <= 65389;
end
4127:begin
x_i <= 65366;
end
4128:begin
x_i <= 65399;
end
4129:begin
x_i <= 65388;
end
4130:begin
x_i <= 65411;
end
4131:begin
x_i <= 65446;
end
4132:begin
x_i <= 65470;
end
4133:begin
x_i <= 65463;
end
4134:begin
x_i <= 65470;
end
4135:begin
x_i <= 65456;
end
4136:begin
x_i <= 65468;
end
4137:begin
x_i <= 65481;
end
4138:begin
x_i <= 65517;
end
4139:begin
x_i <= 65525;
end
4140:begin
x_i <= 17;
end
4141:begin
x_i <= 19;
end
4142:begin
x_i <= 42;
end
4143:begin
x_i <= 65501;
end
4144:begin
x_i <= 20;
end
4145:begin
x_i <= 65527;
end
4146:begin
x_i <= 7;
end
4147:begin
x_i <= 3;
end
4148:begin
x_i <= 65533;
end
4149:begin
x_i <= 38;
end
4150:begin
x_i <= 48;
end
4151:begin
x_i <= 65;
end
4152:begin
x_i <= 107;
end
4153:begin
x_i <= 121;
end
4154:begin
x_i <= 130;
end
4155:begin
x_i <= 99;
end
4156:begin
x_i <= 123;
end
4157:begin
x_i <= 132;
end
4158:begin
x_i <= 135;
end
4159:begin
x_i <= 151;
end
4160:begin
x_i <= 176;
end
4161:begin
x_i <= 123;
end
4162:begin
x_i <= 118;
end
4163:begin
x_i <= 191;
end
4164:begin
x_i <= 235;
end
4165:begin
x_i <= 290;
end
4166:begin
x_i <= 278;
end
4167:begin
x_i <= 384;
end
4168:begin
x_i <= 364;
end
4169:begin
x_i <= 133;
end
4170:begin
x_i <= 5;
end
4171:begin
x_i <= 65402;
end
4172:begin
x_i <= 65341;
end
4173:begin
x_i <= 65292;
end
4174:begin
x_i <= 65287;
end
4175:begin
x_i <= 65425;
end
4176:begin
x_i <= 65427;
end
4177:begin
x_i <= 65433;
end
4178:begin
x_i <= 26;
end
4179:begin
x_i <= 124;
end
4180:begin
x_i <= 66;
end
4181:begin
x_i <= 9;
end
4182:begin
x_i <= 65488;
end
4183:begin
x_i <= 65486;
end
4184:begin
x_i <= 65437;
end
4185:begin
x_i <= 65452;
end
4186:begin
x_i <= 65501;
end
4187:begin
x_i <= 52;
end
4188:begin
x_i <= 21;
end
4189:begin
x_i <= 31;
end
4190:begin
x_i <= 43;
end
4191:begin
x_i <= 38;
end
4192:begin
x_i <= 65495;
end
4193:begin
x_i <= 65420;
end
4194:begin
x_i <= 65391;
end
4195:begin
x_i <= 65426;
end
4196:begin
x_i <= 65433;
end
4197:begin
x_i <= 65507;
end
4198:begin
x_i <= 33;
end
4199:begin
x_i <= 44;
end
4200:begin
x_i <= 10;
end
4201:begin
x_i <= 65515;
end
4202:begin
x_i <= 65489;
end
4203:begin
x_i <= 65396;
end
4204:begin
x_i <= 65343;
end
4205:begin
x_i <= 65292;
end
4206:begin
x_i <= 65326;
end
4207:begin
x_i <= 65379;
end
4208:begin
x_i <= 65454;
end
4209:begin
x_i <= 0;
end
4210:begin
x_i <= 56;
end
4211:begin
x_i <= 65521;
end
4212:begin
x_i <= 65520;
end
4213:begin
x_i <= 12;
end
4214:begin
x_i <= 65475;
end
4215:begin
x_i <= 65423;
end
4216:begin
x_i <= 65426;
end
4217:begin
x_i <= 65389;
end
4218:begin
x_i <= 65391;
end
4219:begin
x_i <= 65338;
end
4220:begin
x_i <= 65327;
end
4221:begin
x_i <= 65364;
end
4222:begin
x_i <= 65353;
end
4223:begin
x_i <= 65380;
end
4224:begin
x_i <= 65340;
end
4225:begin
x_i <= 65379;
end
4226:begin
x_i <= 65406;
end
4227:begin
x_i <= 65371;
end
4228:begin
x_i <= 65401;
end
4229:begin
x_i <= 65401;
end
4230:begin
x_i <= 65340;
end
4231:begin
x_i <= 65339;
end
4232:begin
x_i <= 65354;
end
4233:begin
x_i <= 65383;
end
4234:begin
x_i <= 65391;
end
4235:begin
x_i <= 65408;
end
4236:begin
x_i <= 65431;
end
4237:begin
x_i <= 65447;
end
4238:begin
x_i <= 65469;
end
4239:begin
x_i <= 65463;
end
4240:begin
x_i <= 65484;
end
4241:begin
x_i <= 65483;
end
4242:begin
x_i <= 65463;
end
4243:begin
x_i <= 9;
end
4244:begin
x_i <= 30;
end
4245:begin
x_i <= 13;
end
4246:begin
x_i <= 44;
end
4247:begin
x_i <= 46;
end
4248:begin
x_i <= 46;
end
4249:begin
x_i <= 30;
end
4250:begin
x_i <= 33;
end
4251:begin
x_i <= 8;
end
4252:begin
x_i <= 65504;
end
4253:begin
x_i <= 65505;
end
4254:begin
x_i <= 65526;
end
4255:begin
x_i <= 20;
end
4256:begin
x_i <= 10;
end
4257:begin
x_i <= 90;
end
4258:begin
x_i <= 110;
end
4259:begin
x_i <= 126;
end
4260:begin
x_i <= 130;
end
4261:begin
x_i <= 161;
end
4262:begin
x_i <= 165;
end
4263:begin
x_i <= 142;
end
4264:begin
x_i <= 92;
end
4265:begin
x_i <= 122;
end
4266:begin
x_i <= 163;
end
4267:begin
x_i <= 135;
end
4268:begin
x_i <= 178;
end
4269:begin
x_i <= 156;
end
4270:begin
x_i <= 171;
end
4271:begin
x_i <= 187;
end
4272:begin
x_i <= 182;
end
4273:begin
x_i <= 211;
end
4274:begin
x_i <= 199;
end
4275:begin
x_i <= 210;
end
4276:begin
x_i <= 305;
end
4277:begin
x_i <= 389;
end
4278:begin
x_i <= 282;
end
4279:begin
x_i <= 50;
end
4280:begin
x_i <= 65473;
end
4281:begin
x_i <= 65392;
end
4282:begin
x_i <= 65333;
end
4283:begin
x_i <= 65204;
end
4284:begin
x_i <= 65282;
end
4285:begin
x_i <= 65390;
end
4286:begin
x_i <= 65381;
end
4287:begin
x_i <= 65512;
end
4288:begin
x_i <= 140;
end
4289:begin
x_i <= 163;
end
4290:begin
x_i <= 60;
end
4291:begin
x_i <= 65472;
end
4292:begin
x_i <= 65439;
end
4293:begin
x_i <= 65392;
end
4294:begin
x_i <= 65401;
end
4295:begin
x_i <= 65422;
end
4296:begin
x_i <= 65479;
end
4297:begin
x_i <= 65531;
end
4298:begin
x_i <= 70;
end
4299:begin
x_i <= 40;
end
4300:begin
x_i <= 42;
end
4301:begin
x_i <= 65527;
end
4302:begin
x_i <= 65381;
end
4303:begin
x_i <= 65338;
end
4304:begin
x_i <= 65315;
end
4305:begin
x_i <= 65329;
end
4306:begin
x_i <= 65377;
end
4307:begin
x_i <= 65451;
end
4308:begin
x_i <= 65518;
end
4309:begin
x_i <= 12;
end
4310:begin
x_i <= 65533;
end
4311:begin
x_i <= 65531;
end
4312:begin
x_i <= 65438;
end
4313:begin
x_i <= 65339;
end
4314:begin
x_i <= 65308;
end
4315:begin
x_i <= 65312;
end
4316:begin
x_i <= 65352;
end
4317:begin
x_i <= 65392;
end
4318:begin
x_i <= 65511;
end
4319:begin
x_i <= 48;
end
4320:begin
x_i <= 67;
end
4321:begin
x_i <= 80;
end
4322:begin
x_i <= 38;
end
4323:begin
x_i <= 65495;
end
4324:begin
x_i <= 65438;
end
4325:begin
x_i <= 65438;
end
4326:begin
x_i <= 65392;
end
4327:begin
x_i <= 65433;
end
4328:begin
x_i <= 65401;
end
4329:begin
x_i <= 65443;
end
4330:begin
x_i <= 65478;
end
4331:begin
x_i <= 65477;
end
4332:begin
x_i <= 65495;
end
4333:begin
x_i <= 65495;
end
4334:begin
x_i <= 65450;
end
4335:begin
x_i <= 65441;
end
4336:begin
x_i <= 65372;
end
4337:begin
x_i <= 65367;
end
4338:begin
x_i <= 65449;
end
4339:begin
x_i <= 65404;
end
4340:begin
x_i <= 65457;
end
4341:begin
x_i <= 65469;
end
4342:begin
x_i <= 65429;
end
4343:begin
x_i <= 65435;
end
4344:begin
x_i <= 65396;
end
4345:begin
x_i <= 65367;
end
4346:begin
x_i <= 65368;
end
4347:begin
x_i <= 65371;
end
4348:begin
x_i <= 65370;
end
4349:begin
x_i <= 65461;
end
4350:begin
x_i <= 65484;
end
4351:begin
x_i <= 65530;
end
4352:begin
x_i <= 18;
end
4353:begin
x_i <= 65519;
end
4354:begin
x_i <= 65488;
end
4355:begin
x_i <= 65480;
end
4356:begin
x_i <= 65442;
end
4357:begin
x_i <= 65441;
end
4358:begin
x_i <= 65477;
end
4359:begin
x_i <= 65488;
end
4360:begin
x_i <= 13;
end
4361:begin
x_i <= 3;
end
4362:begin
x_i <= 28;
end
4363:begin
x_i <= 27;
end
4364:begin
x_i <= 4;
end
4365:begin
x_i <= 14;
end
4366:begin
x_i <= 21;
end
4367:begin
x_i <= 14;
end
4368:begin
x_i <= 15;
end
4369:begin
x_i <= 65532;
end
4370:begin
x_i <= 43;
end
4371:begin
x_i <= 78;
end
4372:begin
x_i <= 67;
end
4373:begin
x_i <= 79;
end
4374:begin
x_i <= 46;
end
4375:begin
x_i <= 71;
end
4376:begin
x_i <= 38;
end
4377:begin
x_i <= 28;
end
4378:begin
x_i <= 68;
end
4379:begin
x_i <= 94;
end
4380:begin
x_i <= 121;
end
4381:begin
x_i <= 124;
end
4382:begin
x_i <= 161;
end
4383:begin
x_i <= 175;
end
4384:begin
x_i <= 135;
end
4385:begin
x_i <= 147;
end
4386:begin
x_i <= 153;
end
4387:begin
x_i <= 174;
end
4388:begin
x_i <= 190;
end
4389:begin
x_i <= 204;
end
4390:begin
x_i <= 218;
end
4391:begin
x_i <= 245;
end
4392:begin
x_i <= 226;
end
4393:begin
x_i <= 154;
end
4394:begin
x_i <= 27;
end
4395:begin
x_i <= 65451;
end
4396:begin
x_i <= 65399;
end
4397:begin
x_i <= 65334;
end
4398:begin
x_i <= 65359;
end
4399:begin
x_i <= 65402;
end
4400:begin
x_i <= 65506;
end
4401:begin
x_i <= 12;
end
4402:begin
x_i <= 61;
end
4403:begin
x_i <= 90;
end
4404:begin
x_i <= 47;
end
4405:begin
x_i <= 4;
end
4406:begin
x_i <= 65467;
end
4407:begin
x_i <= 65471;
end
4408:begin
x_i <= 65452;
end
4409:begin
x_i <= 65445;
end
4410:begin
x_i <= 65496;
end
4411:begin
x_i <= 21;
end
4412:begin
x_i <= 13;
end
4413:begin
x_i <= 39;
end
4414:begin
x_i <= 33;
end
4415:begin
x_i <= 65535;
end
4416:begin
x_i <= 65489;
end
4417:begin
x_i <= 65432;
end
4418:begin
x_i <= 65415;
end
4419:begin
x_i <= 65436;
end
4420:begin
x_i <= 65464;
end
4421:begin
x_i <= 65509;
end
4422:begin
x_i <= 65529;
end
4423:begin
x_i <= 23;
end
4424:begin
x_i <= 28;
end
4425:begin
x_i <= 65528;
end
4426:begin
x_i <= 65468;
end
4427:begin
x_i <= 65424;
end
4428:begin
x_i <= 65386;
end
4429:begin
x_i <= 65358;
end
4430:begin
x_i <= 65391;
end
4431:begin
x_i <= 65423;
end
4432:begin
x_i <= 65453;
end
4433:begin
x_i <= 65524;
end
4434:begin
x_i <= 27;
end
4435:begin
x_i <= 36;
end
4436:begin
x_i <= 1;
end
4437:begin
x_i <= 65487;
end
4438:begin
x_i <= 65448;
end
4439:begin
x_i <= 65441;
end
4440:begin
x_i <= 65447;
end
4441:begin
x_i <= 65422;
end
4442:begin
x_i <= 65465;
end
4443:begin
x_i <= 65474;
end
4444:begin
x_i <= 65466;
end
4445:begin
x_i <= 65447;
end
4446:begin
x_i <= 65431;
end
4447:begin
x_i <= 65451;
end
4448:begin
x_i <= 65416;
end
4449:begin
x_i <= 65409;
end
4450:begin
x_i <= 65436;
end
4451:begin
x_i <= 65466;
end
4452:begin
x_i <= 65457;
end
4453:begin
x_i <= 65441;
end
4454:begin
x_i <= 65453;
end
4455:begin
x_i <= 65454;
end
4456:begin
x_i <= 65434;
end
4457:begin
x_i <= 65481;
end
4458:begin
x_i <= 65405;
end
4459:begin
x_i <= 65392;
end
4460:begin
x_i <= 65370;
end
4461:begin
x_i <= 65366;
end
4462:begin
x_i <= 65392;
end
4463:begin
x_i <= 65402;
end
4464:begin
x_i <= 65393;
end
4465:begin
x_i <= 65410;
end
4466:begin
x_i <= 65441;
end
4467:begin
x_i <= 65404;
end
4468:begin
x_i <= 65431;
end
4469:begin
x_i <= 65423;
end
4470:begin
x_i <= 65410;
end
4471:begin
x_i <= 65429;
end
4472:begin
x_i <= 65406;
end
4473:begin
x_i <= 65482;
end
4474:begin
x_i <= 1;
end
4475:begin
x_i <= 65533;
end
4476:begin
x_i <= 16;
end
4477:begin
x_i <= 52;
end
4478:begin
x_i <= 30;
end
4479:begin
x_i <= 19;
end
4480:begin
x_i <= 65508;
end
4481:begin
x_i <= 65497;
end
4482:begin
x_i <= 17;
end
4483:begin
x_i <= 35;
end
4484:begin
x_i <= 44;
end
4485:begin
x_i <= 87;
end
4486:begin
x_i <= 96;
end
4487:begin
x_i <= 107;
end
4488:begin
x_i <= 89;
end
4489:begin
x_i <= 84;
end
4490:begin
x_i <= 59;
end
4491:begin
x_i <= 56;
end
4492:begin
x_i <= 43;
end
4493:begin
x_i <= 65;
end
4494:begin
x_i <= 36;
end
4495:begin
x_i <= 46;
end
4496:begin
x_i <= 71;
end
4497:begin
x_i <= 97;
end
4498:begin
x_i <= 129;
end
4499:begin
x_i <= 113;
end
4500:begin
x_i <= 110;
end
4501:begin
x_i <= 71;
end
4502:begin
x_i <= 94;
end
4503:begin
x_i <= 69;
end
4504:begin
x_i <= 49;
end
4505:begin
x_i <= 99;
end
4506:begin
x_i <= 89;
end
4507:begin
x_i <= 102;
end
4508:begin
x_i <= 118;
end
4509:begin
x_i <= 102;
end
4510:begin
x_i <= 139;
end
4511:begin
x_i <= 145;
end
4512:begin
x_i <= 121;
end
4513:begin
x_i <= 147;
end
4514:begin
x_i <= 126;
end
4515:begin
x_i <= 99;
end
4516:begin
x_i <= 86;
end
4517:begin
x_i <= 78;
end
4518:begin
x_i <= 44;
end
4519:begin
x_i <= 33;
end
4520:begin
x_i <= 65502;
end
4521:begin
x_i <= 65455;
end
4522:begin
x_i <= 65448;
end
4523:begin
x_i <= 65428;
end
4524:begin
x_i <= 65465;
end
4525:begin
x_i <= 65480;
end
4526:begin
x_i <= 65486;
end
4527:begin
x_i <= 65486;
end
4528:begin
x_i <= 65488;
end
4529:begin
x_i <= 65493;
end
4530:begin
x_i <= 65483;
end
4531:begin
x_i <= 65457;
end
4532:begin
x_i <= 65487;
end
4533:begin
x_i <= 65454;
end
4534:begin
x_i <= 65498;
end
4535:begin
x_i <= 65491;
end
4536:begin
x_i <= 65499;
end
4537:begin
x_i <= 65512;
end
4538:begin
x_i <= 65504;
end
4539:begin
x_i <= 65487;
end
4540:begin
x_i <= 65486;
end
4541:begin
x_i <= 65470;
end
4542:begin
x_i <= 65431;
end
4543:begin
x_i <= 65421;
end
4544:begin
x_i <= 65422;
end
4545:begin
x_i <= 65460;
end
4546:begin
x_i <= 65450;
end
4547:begin
x_i <= 65436;
end
4548:begin
x_i <= 65442;
end
4549:begin
x_i <= 65452;
end
4550:begin
x_i <= 65466;
end
4551:begin
x_i <= 65460;
end
4552:begin
x_i <= 65456;
end
4553:begin
x_i <= 65448;
end
4554:begin
x_i <= 65415;
end
4555:begin
x_i <= 65427;
end
4556:begin
x_i <= 65426;
end
4557:begin
x_i <= 65462;
end
4558:begin
x_i <= 65463;
end
4559:begin
x_i <= 65479;
end
4560:begin
x_i <= 65488;
end
4561:begin
x_i <= 65511;
end
4562:begin
x_i <= 65496;
end
4563:begin
x_i <= 65459;
end
4564:begin
x_i <= 65441;
end
4565:begin
x_i <= 65421;
end
4566:begin
x_i <= 65437;
end
4567:begin
x_i <= 65460;
end
4568:begin
x_i <= 65456;
end
4569:begin
x_i <= 65470;
end
4570:begin
x_i <= 65485;
end
4571:begin
x_i <= 65500;
end
4572:begin
x_i <= 65504;
end
4573:begin
x_i <= 65456;
end
4574:begin
x_i <= 65499;
end
4575:begin
x_i <= 65492;
end
4576:begin
x_i <= 65480;
end
4577:begin
x_i <= 65496;
end
4578:begin
x_i <= 65507;
end
4579:begin
x_i <= 65469;
end
4580:begin
x_i <= 65472;
end
4581:begin
x_i <= 65407;
end
4582:begin
x_i <= 65436;
end
4583:begin
x_i <= 65401;
end
4584:begin
x_i <= 65394;
end
4585:begin
x_i <= 65429;
end
4586:begin
x_i <= 65444;
end
4587:begin
x_i <= 65494;
end
4588:begin
x_i <= 12;
end
4589:begin
x_i <= 65461;
end
4590:begin
x_i <= 65522;
end
4591:begin
x_i <= 65474;
end
4592:begin
x_i <= 65500;
end
4593:begin
x_i <= 65527;
end
4594:begin
x_i <= 65482;
end
4595:begin
x_i <= 65527;
end
4596:begin
x_i <= 65522;
end
4597:begin
x_i <= 65493;
end
4598:begin
x_i <= 65507;
end
4599:begin
x_i <= 65511;
end
4600:begin
x_i <= 65515;
end
4601:begin
x_i <= 65508;
end
4602:begin
x_i <= 65513;
end
4603:begin
x_i <= 65527;
end
4604:begin
x_i <= 11;
end
4605:begin
x_i <= 65535;
end
4606:begin
x_i <= 5;
end
4607:begin
x_i <= 57;
end
4608:begin
x_i <= 61;
end
4609:begin
x_i <= 101;
end
4610:begin
x_i <= 40;
end
4611:begin
x_i <= 68;
end
4612:begin
x_i <= 89;
end
4613:begin
x_i <= 30;
end
4614:begin
x_i <= 36;
end
4615:begin
x_i <= 11;
end
4616:begin
x_i <= 10;
end
4617:begin
x_i <= 65514;
end
4618:begin
x_i <= 11;
end
4619:begin
x_i <= 65;
end
4620:begin
x_i <= 101;
end
4621:begin
x_i <= 91;
end
4622:begin
x_i <= 99;
end
4623:begin
x_i <= 98;
end
4624:begin
x_i <= 72;
end
4625:begin
x_i <= 78;
end
4626:begin
x_i <= 71;
end
4627:begin
x_i <= 91;
end
4628:begin
x_i <= 90;
end
4629:begin
x_i <= 98;
end
4630:begin
x_i <= 80;
end
4631:begin
x_i <= 79;
end
4632:begin
x_i <= 88;
end
4633:begin
x_i <= 74;
end
4634:begin
x_i <= 107;
end
4635:begin
x_i <= 98;
end
4636:begin
x_i <= 128;
end
4637:begin
x_i <= 186;
end
4638:begin
x_i <= 165;
end
4639:begin
x_i <= 129;
end
4640:begin
x_i <= 94;
end
4641:begin
x_i <= 5;
end
4642:begin
x_i <= 65457;
end
4643:begin
x_i <= 65351;
end
4644:begin
x_i <= 65368;
end
4645:begin
x_i <= 65351;
end
4646:begin
x_i <= 65363;
end
4647:begin
x_i <= 65443;
end
4648:begin
x_i <= 65496;
end
4649:begin
x_i <= 65521;
end
4650:begin
x_i <= 65531;
end
4651:begin
x_i <= 65500;
end
4652:begin
x_i <= 65507;
end
4653:begin
x_i <= 65469;
end
4654:begin
x_i <= 65416;
end
4655:begin
x_i <= 65452;
end
4656:begin
x_i <= 65486;
end
4657:begin
x_i <= 65483;
end
4658:begin
x_i <= 65506;
end
4659:begin
x_i <= 10;
end
4660:begin
x_i <= 65528;
end
4661:begin
x_i <= 65523;
end
4662:begin
x_i <= 65476;
end
4663:begin
x_i <= 65458;
end
4664:begin
x_i <= 65439;
end
4665:begin
x_i <= 65417;
end
4666:begin
x_i <= 65437;
end
4667:begin
x_i <= 65489;
end
4668:begin
x_i <= 65471;
end
4669:begin
x_i <= 65502;
end
4670:begin
x_i <= 65529;
end
4671:begin
x_i <= 65482;
end
4672:begin
x_i <= 65509;
end
4673:begin
x_i <= 65510;
end
4674:begin
x_i <= 65462;
end
4675:begin
x_i <= 65442;
end
4676:begin
x_i <= 65441;
end
4677:begin
x_i <= 65438;
end
4678:begin
x_i <= 65445;
end
4679:begin
x_i <= 65455;
end
4680:begin
x_i <= 65526;
end
4681:begin
x_i <= 20;
end
4682:begin
x_i <= 9;
end
4683:begin
x_i <= 23;
end
4684:begin
x_i <= 65531;
end
4685:begin
x_i <= 16;
end
4686:begin
x_i <= 5;
end
4687:begin
x_i <= 65518;
end
4688:begin
x_i <= 65481;
end
4689:begin
x_i <= 65472;
end
4690:begin
x_i <= 65520;
end
4691:begin
x_i <= 65498;
end
4692:begin
x_i <= 65497;
end
4693:begin
x_i <= 4;
end
4694:begin
x_i <= 24;
end
4695:begin
x_i <= 18;
end
4696:begin
x_i <= 21;
end
4697:begin
x_i <= 65531;
end
4698:begin
x_i <= 47;
end
4699:begin
x_i <= 65535;
end
4700:begin
x_i <= 65531;
end
4701:begin
x_i <= 65535;
end
4702:begin
x_i <= 65531;
end
4703:begin
x_i <= 65527;
end
4704:begin
x_i <= 65534;
end
4705:begin
x_i <= 65503;
end
4706:begin
x_i <= 65511;
end
4707:begin
x_i <= 65429;
end
4708:begin
x_i <= 65353;
end
4709:begin
x_i <= 65363;
end
4710:begin
x_i <= 65319;
end
4711:begin
x_i <= 65371;
end
4712:begin
x_i <= 65391;
end
4713:begin
x_i <= 65443;
end
4714:begin
x_i <= 5;
end
4715:begin
x_i <= 65510;
end
4716:begin
x_i <= 65531;
end
4717:begin
x_i <= 65523;
end
4718:begin
x_i <= 65472;
end
4719:begin
x_i <= 65430;
end
4720:begin
x_i <= 65393;
end
4721:begin
x_i <= 65364;
end
4722:begin
x_i <= 65417;
end
4723:begin
x_i <= 65402;
end
4724:begin
x_i <= 65428;
end
4725:begin
x_i <= 65507;
end
4726:begin
x_i <= 65492;
end
4727:begin
x_i <= 65517;
end
4728:begin
x_i <= 65523;
end
4729:begin
x_i <= 65478;
end
4730:begin
x_i <= 65444;
end
4731:begin
x_i <= 65442;
end
4732:begin
x_i <= 65427;
end
4733:begin
x_i <= 65491;
end
4734:begin
x_i <= 12;
end
4735:begin
x_i <= 1;
end
4736:begin
x_i <= 66;
end
4737:begin
x_i <= 42;
end
4738:begin
x_i <= 36;
end
4739:begin
x_i <= 5;
end
4740:begin
x_i <= 65490;
end
4741:begin
x_i <= 65492;
end
4742:begin
x_i <= 65493;
end
4743:begin
x_i <= 65470;
end
4744:begin
x_i <= 39;
end
4745:begin
x_i <= 61;
end
4746:begin
x_i <= 71;
end
4747:begin
x_i <= 99;
end
4748:begin
x_i <= 125;
end
4749:begin
x_i <= 92;
end
4750:begin
x_i <= 82;
end
4751:begin
x_i <= 86;
end
4752:begin
x_i <= 23;
end
4753:begin
x_i <= 27;
end
4754:begin
x_i <= 59;
end
4755:begin
x_i <= 30;
end
4756:begin
x_i <= 84;
end
4757:begin
x_i <= 75;
end
4758:begin
x_i <= 134;
end
4759:begin
x_i <= 202;
end
4760:begin
x_i <= 173;
end
4761:begin
x_i <= 193;
end
4762:begin
x_i <= 191;
end
4763:begin
x_i <= 137;
end
4764:begin
x_i <= 52;
end
4765:begin
x_i <= 65483;
end
4766:begin
x_i <= 65354;
end
4767:begin
x_i <= 65349;
end
4768:begin
x_i <= 65343;
end
4769:begin
x_i <= 65338;
end
4770:begin
x_i <= 65418;
end
4771:begin
x_i <= 65505;
end
4772:begin
x_i <= 7;
end
4773:begin
x_i <= 55;
end
4774:begin
x_i <= 45;
end
4775:begin
x_i <= 29;
end
4776:begin
x_i <= 65512;
end
4777:begin
x_i <= 65433;
end
4778:begin
x_i <= 65431;
end
4779:begin
x_i <= 65455;
end
4780:begin
x_i <= 65480;
end
4781:begin
x_i <= 65503;
end
4782:begin
x_i <= 32;
end
4783:begin
x_i <= 60;
end
4784:begin
x_i <= 57;
end
4785:begin
x_i <= 36;
end
4786:begin
x_i <= 65509;
end
4787:begin
x_i <= 65460;
end
4788:begin
x_i <= 65419;
end
4789:begin
x_i <= 65404;
end
4790:begin
x_i <= 65437;
end
4791:begin
x_i <= 65478;
end
4792:begin
x_i <= 65474;
end
4793:begin
x_i <= 20;
end
4794:begin
x_i <= 79;
end
4795:begin
x_i <= 63;
end
4796:begin
x_i <= 72;
end
4797:begin
x_i <= 18;
end
4798:begin
x_i <= 65490;
end
4799:begin
x_i <= 65448;
end
4800:begin
x_i <= 65428;
end
4801:begin
x_i <= 65391;
end
4802:begin
x_i <= 65444;
end
4803:begin
x_i <= 65500;
end
4804:begin
x_i <= 16;
end
4805:begin
x_i <= 55;
end
4806:begin
x_i <= 59;
end
4807:begin
x_i <= 44;
end
4808:begin
x_i <= 1;
end
4809:begin
x_i <= 65506;
end
4810:begin
x_i <= 65489;
end
4811:begin
x_i <= 65442;
end
4812:begin
x_i <= 65428;
end
4813:begin
x_i <= 65430;
end
4814:begin
x_i <= 65488;
end
4815:begin
x_i <= 65480;
end
4816:begin
x_i <= 65499;
end
4817:begin
x_i <= 65520;
end
4818:begin
x_i <= 65513;
end
4819:begin
x_i <= 5;
end
4820:begin
x_i <= 65510;
end
4821:begin
x_i <= 65479;
end
4822:begin
x_i <= 65459;
end
4823:begin
x_i <= 65462;
end
4824:begin
x_i <= 65454;
end
4825:begin
x_i <= 65488;
end
4826:begin
x_i <= 65489;
end
4827:begin
x_i <= 65525;
end
4828:begin
x_i <= 5;
end
4829:begin
x_i <= 65512;
end
4830:begin
x_i <= 65516;
end
4831:begin
x_i <= 65481;
end
4832:begin
x_i <= 65458;
end
4833:begin
x_i <= 65456;
end
4834:begin
x_i <= 65453;
end
4835:begin
x_i <= 65468;
end
4836:begin
x_i <= 65421;
end
4837:begin
x_i <= 65372;
end
4838:begin
x_i <= 65367;
end
4839:begin
x_i <= 65331;
end
4840:begin
x_i <= 65383;
end
4841:begin
x_i <= 65413;
end
4842:begin
x_i <= 65364;
end
4843:begin
x_i <= 65454;
end
4844:begin
x_i <= 65460;
end
4845:begin
x_i <= 65439;
end
4846:begin
x_i <= 65505;
end
4847:begin
x_i <= 65472;
end
4848:begin
x_i <= 65428;
end
4849:begin
x_i <= 65459;
end
4850:begin
x_i <= 65406;
end
4851:begin
x_i <= 65420;
end
4852:begin
x_i <= 65422;
end
4853:begin
x_i <= 65440;
end
4854:begin
x_i <= 65464;
end
4855:begin
x_i <= 65500;
end
4856:begin
x_i <= 65481;
end
4857:begin
x_i <= 65485;
end
4858:begin
x_i <= 65432;
end
4859:begin
x_i <= 65463;
end
4860:begin
x_i <= 65490;
end
4861:begin
x_i <= 65464;
end
4862:begin
x_i <= 65498;
end
4863:begin
x_i <= 5;
end
4864:begin
x_i <= 65514;
end
4865:begin
x_i <= 1;
end
4866:begin
x_i <= 27;
end
4867:begin
x_i <= 26;
end
4868:begin
x_i <= 45;
end
4869:begin
x_i <= 33;
end
4870:begin
x_i <= 65528;
end
4871:begin
x_i <= 65521;
end
4872:begin
x_i <= 65507;
end
4873:begin
x_i <= 65525;
end
4874:begin
x_i <= 11;
end
4875:begin
x_i <= 5;
end
4876:begin
x_i <= 67;
end
4877:begin
x_i <= 120;
end
4878:begin
x_i <= 119;
end
4879:begin
x_i <= 162;
end
4880:begin
x_i <= 0;
end
endcase
end

always begin
	#10
	if(index2==50)begin
			write <= 1;
			index2 <= 0;
		end
		else begin
			index2 <= index2+1;
			write <= 0;
		end
end


always begin
	#500
	if(index==4880)begin
		index <= 0;
	end
	else begin
		index <= index+1;
	end
end
	

	initial begin
		// Initialize Inputs
		clk = 0;
		x_i = 0;
		write = 0;
		reset = 0;
		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

