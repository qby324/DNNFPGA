
 
 
 




window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"


      waveform add -signals /nnpara8bit_tb/status
      waveform add -signals /nnpara8bit_tb/nnpara8bit_synth_inst/bmg_port/CLKA
      waveform add -signals /nnpara8bit_tb/nnpara8bit_synth_inst/bmg_port/ADDRA
      waveform add -signals /nnpara8bit_tb/nnpara8bit_synth_inst/bmg_port/DOUTA
console submit -using simulator -wait no "run"
