`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:05:47 12/16/2011 
// Design Name: 
// Module Name:    log2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//	����:64bit
//	�o��:signed 21bit
//	�ΐ��̐�����:63~0 10000�{
//      �ŏ���bit��1�ɂȂ����ꏊ���ΐ���̐������Ɉ�v����
//	�������̌��10bit���`�F�b�N���đΐ��ɋߎ�
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module log2_10bit(clk,start,indata,outdata,dv);
   input clk;                    //!< Global Clock
   input start;                  //!< module start (active high)
   input [63:0] indata;          //!< InputData  (    X    )
   output signed [20:0] outdata; //!< OutputData ( log2(X) )
   output 		dv;      //!< Data Valid (active high)
   reg 			dv=0;
   reg signed [20:0] 	outdata=0;	
   
   /* Other Register */
   reg [6:0] 		inte=63;    //!< �ΐ��������̐���
   reg [9:0] 		intemp=0;   //!< ����bit�̎������bit
   reg signed [13:0] 	fraction=0; //!< ��������
   reg [2:0] 		clk_cnt=0;  //!< Calclation Process
                                    //!< (0:getdata 1:integer 2:fraction1 3:frac2 4:output)
   reg [6:0] 		i=63;
   
   always@(posedge clk) begin
      if(start==1) begin	//!< Start Log Calculation

	 /*  Calc Integer  */
	 if(inte==0)begin
	    dv<=1;
	    outdata<=0;
	 end else begin
	    
	    case(clk_cnt)
	      0:begin
		 if(indata[63:50]==14'b0)begin
		    inte<=49;
		 end else if(indata[49:40]==10'b0)begin
		    inte<=39;
		 end else begin
		    inte<=63;
		 end
		 clk_cnt<=1;
	      end
	      1:begin
		 if(indata[inte]==1)begin
		    clk_cnt<=2;
		 end else begin
		    inte<=inte-1;
		 end
	      end
	      2:begin
		 clk_cnt<=3;
		 /* Calc fraction          */
		 /* 1�ɂȂ���bit�ʒu�̐^����10bit���������Z */
		 /* �����̈ʒu�ɂ���Ă��낢��ς��� */
		 if(inte>=10)
		   intemp<={indata[inte-1],indata[inte-2],indata[inte-3],indata[inte-4],indata[inte-5],indata[inte-6],indata[inte-7],indata[inte-8],indata[inte-9],indata[inte-10]};
		 else if(inte==9)
		   intemp<={indata[inte-1],indata[inte-2],indata[inte-3],indata[inte-4],indata[inte-5],indata[inte-6],indata[inte-7],indata[inte-8],indata[inte-9],1'b0};
		 else if(inte==8)
		   intemp<={indata[inte-1],indata[inte-2],indata[inte-3],indata[inte-4],indata[inte-5],indata[inte-6],indata[inte-7],indata[inte-8],2'b0};
		 else if(inte==7)
		   intemp<={indata[inte-1],indata[inte-2],indata[inte-3],indata[inte-4],indata[inte-5],indata[inte-6],indata[inte-7],3'b0};
		 else if(inte==6)
		   intemp<={indata[inte-1],indata[inte-2],indata[inte-3],indata[inte-4],indata[inte-5],indata[inte-6],4'b0};
		 else if(inte==5)
		   intemp<={indata[inte-1],indata[inte-2],indata[inte-3],indata[inte-4],indata[inte-5],5'b0};
		 else if(inte==4)
		   intemp<={indata[inte-1],indata[inte-2],indata[inte-3],indata[inte-4],6'b0};
		 else if(inte==3)
		   intemp<={indata[inte-1],indata[inte-2],indata[inte-3],7'b0};
		 else if(inte==2)
		   intemp<={indata[inte-1],indata[inte-2],8'b0};
		 else if(inte==1)
		   intemp<={indata[inte-1],9'b0};
		 else if(inte==0)
		   intemp<=10'b0;
	      end
	      3:begin
		 clk_cnt<=4;
		 //�����̃e�[�u��
		 case(intemp)
		0	:fraction <= 0;
		1	:fraction <= 23;
		2	:fraction <= 46;
		3	:fraction <= 69;
		4	:fraction <= 92;
		5	:fraction <= 115;
		6	:fraction <= 138;
		7	:fraction <= 161;
		8	:fraction <= 183;
		9	:fraction <= 206;
		10	:fraction <= 229;
		11	:fraction <= 252;
		12	:fraction <= 275;
		13	:fraction <= 298;
		14	:fraction <= 320;
		15	:fraction <= 343;
		16	:fraction <= 366;
		17	:fraction <= 389;
		18	:fraction <= 411;
		19	:fraction <= 434;
		20	:fraction <= 457;
		21	:fraction <= 479;
		22	:fraction <= 502;
		23	:fraction <= 525;
		24	:fraction <= 547;
		25	:fraction <= 570;
		26	:fraction <= 592;
		27	:fraction <= 615;
		28	:fraction <= 637;
		29	:fraction <= 660;
		30	:fraction <= 682;
		31	:fraction <= 704;
		32	:fraction <= 727;
		33	:fraction <= 749;
		34	:fraction <= 772;
		35	:fraction <= 794;
		36	:fraction <= 816;
		37	:fraction <= 839;
		38	:fraction <= 861;
		39	:fraction <= 883;
		40	:fraction <= 905;
		41	:fraction <= 927;
		42	:fraction <= 950;
		43	:fraction <= 972;
		44	:fraction <= 994;
		45	:fraction <= 1016;
		46	:fraction <= 1038;
		47	:fraction <= 1060;
		48	:fraction <= 1082;
		49	:fraction <= 1104;
		50	:fraction <= 1126;
		51	:fraction <= 1148;
		52	:fraction <= 1170;
		53	:fraction <= 1192;
		54	:fraction <= 1214;
		55	:fraction <= 1236;
		56	:fraction <= 1258;
		57	:fraction <= 1280;
		58	:fraction <= 1302;
		59	:fraction <= 1324;
		60	:fraction <= 1345;
		61	:fraction <= 1367;
		62	:fraction <= 1389;
		63	:fraction <= 1411;
		64	:fraction <= 1432;
		65	:fraction <= 1454;
		66	:fraction <= 1476;
		67	:fraction <= 1498;
		68	:fraction <= 1519;
		69	:fraction <= 1541;
		70	:fraction <= 1562;
		71	:fraction <= 1584;
		72	:fraction <= 1606;
		73	:fraction <= 1627;
		74	:fraction <= 1649;
		75	:fraction <= 1670;
		76	:fraction <= 1692;
		77	:fraction <= 1713;
		78	:fraction <= 1735;
		79	:fraction <= 1756;
		80	:fraction <= 1778;
		81	:fraction <= 1799;
		82	:fraction <= 1820;
		83	:fraction <= 1842;
		84	:fraction <= 1863;
		85	:fraction <= 1884;
		86	:fraction <= 1906;
		87	:fraction <= 1927;
		88	:fraction <= 1948;
		89	:fraction <= 1969;
		90	:fraction <= 1991;
		91	:fraction <= 2012;
		92	:fraction <= 2033;
		93	:fraction <= 2054;
		94	:fraction <= 2075;
		95	:fraction <= 2097;
		96	:fraction <= 2118;
		97	:fraction <= 2139;
		98	:fraction <= 2160;
		99	:fraction <= 2181;
		100	:fraction <= 2202;
		101	:fraction <= 2223;
		102	:fraction <= 2244;
		103	:fraction <= 2265;
		104	:fraction <= 2286;
		105	:fraction <= 2307;
		106	:fraction <= 2328;
		107	:fraction <= 2349;
		108	:fraction <= 2370;
		109	:fraction <= 2390;
		110	:fraction <= 2411;
		111	:fraction <= 2432;
		112	:fraction <= 2453;
		113	:fraction <= 2474;
		114	:fraction <= 2495;
		115	:fraction <= 2515;
		116	:fraction <= 2536;
		117	:fraction <= 2557;
		118	:fraction <= 2577;
		119	:fraction <= 2598;
		120	:fraction <= 2619;
		121	:fraction <= 2639;
		122	:fraction <= 2660;
		123	:fraction <= 2681;
		124	:fraction <= 2701;
		125	:fraction <= 2722;
		126	:fraction <= 2742;
		127	:fraction <= 2763;
		128	:fraction <= 2784;
		129	:fraction <= 2804;
		130	:fraction <= 2825;
		131	:fraction <= 2845;
		132	:fraction <= 2865;
		133	:fraction <= 2886;
		134	:fraction <= 2906;
		135	:fraction <= 2927;
		136	:fraction <= 2947;
		137	:fraction <= 2967;
		138	:fraction <= 2988;
		139	:fraction <= 3008;
		140	:fraction <= 3028;
		141	:fraction <= 3049;
		142	:fraction <= 3069;
		143	:fraction <= 3089;
		144	:fraction <= 3110;
		145	:fraction <= 3130;
		146	:fraction <= 3150;
		147	:fraction <= 3170;
		148	:fraction <= 3190;
		149	:fraction <= 3211;
		150	:fraction <= 3231;
		151	:fraction <= 3251;
		152	:fraction <= 3271;
		153	:fraction <= 3291;
		154	:fraction <= 3311;
		155	:fraction <= 3331;
		156	:fraction <= 3351;
		157	:fraction <= 3371;
		158	:fraction <= 3391;
		159	:fraction <= 3411;
		160	:fraction <= 3431;
		161	:fraction <= 3451;
		162	:fraction <= 3471;
		163	:fraction <= 3491;
		164	:fraction <= 3511;
		165	:fraction <= 3531;
		166	:fraction <= 3551;
		167	:fraction <= 3571;
		168	:fraction <= 3590;
		169	:fraction <= 3610;
		170	:fraction <= 3630;
		171	:fraction <= 3650;
		172	:fraction <= 3670;
		173	:fraction <= 3689;
		174	:fraction <= 3709;
		175	:fraction <= 3729;
		176	:fraction <= 3748;
		177	:fraction <= 3768;
		178	:fraction <= 3788;
		179	:fraction <= 3807;
		180	:fraction <= 3827;
		181	:fraction <= 3847;
		182	:fraction <= 3866;
		183	:fraction <= 3886;
		184	:fraction <= 3906;
		185	:fraction <= 3925;
		186	:fraction <= 3945;
		187	:fraction <= 3964;
		188	:fraction <= 3984;
		189	:fraction <= 4003;
		190	:fraction <= 4023;
		191	:fraction <= 4042;
		192	:fraction <= 4062;
		193	:fraction <= 4081;
		194	:fraction <= 4100;
		195	:fraction <= 4120;
		196	:fraction <= 4139;
		197	:fraction <= 4159;
		198	:fraction <= 4178;
		199	:fraction <= 4197;
		200	:fraction <= 4217;
		201	:fraction <= 4236;
		202	:fraction <= 4255;
		203	:fraction <= 4274;
		204	:fraction <= 4294;
		205	:fraction <= 4313;
		206	:fraction <= 4332;
		207	:fraction <= 4351;
		208	:fraction <= 4371;
		209	:fraction <= 4390;
		210	:fraction <= 4409;
		211	:fraction <= 4428;
		212	:fraction <= 4447;
		213	:fraction <= 4466;
		214	:fraction <= 4485;
		215	:fraction <= 4504;
		216	:fraction <= 4524;
		217	:fraction <= 4543;
		218	:fraction <= 4562;
		219	:fraction <= 4581;
		220	:fraction <= 4600;
		221	:fraction <= 4619;
		222	:fraction <= 4638;
		223	:fraction <= 4657;
		224	:fraction <= 4676;
		225	:fraction <= 4694;
		226	:fraction <= 4713;
		227	:fraction <= 4732;
		228	:fraction <= 4751;
		229	:fraction <= 4770;
		230	:fraction <= 4789;
		231	:fraction <= 4808;
		232	:fraction <= 4827;
		233	:fraction <= 4845;
		234	:fraction <= 4864;
		235	:fraction <= 4883;
		236	:fraction <= 4902;
		237	:fraction <= 4920;
		238	:fraction <= 4939;
		239	:fraction <= 4958;
		240	:fraction <= 4977;
		241	:fraction <= 4995;
		242	:fraction <= 5014;
		243	:fraction <= 5033;
		244	:fraction <= 5051;
		245	:fraction <= 5070;
		246	:fraction <= 5089;
		247	:fraction <= 5107;
		248	:fraction <= 5126;
		249	:fraction <= 5144;
		250	:fraction <= 5163;
		251	:fraction <= 5181;
		252	:fraction <= 5200;
		253	:fraction <= 5219;
		254	:fraction <= 5237;
		255	:fraction <= 5255;
		256	:fraction <= 5274;
		257	:fraction <= 5292;
		258	:fraction <= 5311;
		259	:fraction <= 5329;
		260	:fraction <= 5348;
		261	:fraction <= 5366;
		262	:fraction <= 5385;
		263	:fraction <= 5403;
		264	:fraction <= 5421;
		265	:fraction <= 5440;
		266	:fraction <= 5458;
		267	:fraction <= 5476;
		268	:fraction <= 5495;
		269	:fraction <= 5513;
		270	:fraction <= 5531;
		271	:fraction <= 5549;
		272	:fraction <= 5568;
		273	:fraction <= 5586;
		274	:fraction <= 5604;
		275	:fraction <= 5622;
		276	:fraction <= 5640;
		277	:fraction <= 5659;
		278	:fraction <= 5677;
		279	:fraction <= 5695;
		280	:fraction <= 5713;
		281	:fraction <= 5731;
		282	:fraction <= 5749;
		283	:fraction <= 5767;
		284	:fraction <= 5785;
		285	:fraction <= 5804;
		286	:fraction <= 5822;
		287	:fraction <= 5840;
		288	:fraction <= 5858;
		289	:fraction <= 5876;
		290	:fraction <= 5894;
		291	:fraction <= 5912;
		292	:fraction <= 5930;
		293	:fraction <= 5948;
		294	:fraction <= 5965;
		295	:fraction <= 5983;
		296	:fraction <= 6001;
		297	:fraction <= 6019;
		298	:fraction <= 6037;
		299	:fraction <= 6055;
		300	:fraction <= 6073;
		301	:fraction <= 6091;
		302	:fraction <= 6109;
		303	:fraction <= 6126;
		304	:fraction <= 6144;
		305	:fraction <= 6162;
		306	:fraction <= 6180;
		307	:fraction <= 6197;
		308	:fraction <= 6215;
		309	:fraction <= 6233;
		310	:fraction <= 6251;
		311	:fraction <= 6268;
		312	:fraction <= 6286;
		313	:fraction <= 6304;
		314	:fraction <= 6321;
		315	:fraction <= 6339;
		316	:fraction <= 6357;
		317	:fraction <= 6374;
		318	:fraction <= 6392;
		319	:fraction <= 6410;
		320	:fraction <= 6427;
		321	:fraction <= 6445;
		322	:fraction <= 6462;
		323	:fraction <= 6480;
		324	:fraction <= 6497;
		325	:fraction <= 6515;
		326	:fraction <= 6533;
		327	:fraction <= 6550;
		328	:fraction <= 6568;
		329	:fraction <= 6585;
		330	:fraction <= 6602;
		331	:fraction <= 6620;
		332	:fraction <= 6637;
		333	:fraction <= 6655;
		334	:fraction <= 6672;
		335	:fraction <= 6690;
		336	:fraction <= 6707;
		337	:fraction <= 6724;
		338	:fraction <= 6742;
		339	:fraction <= 6759;
		340	:fraction <= 6776;
		341	:fraction <= 6794;
		342	:fraction <= 6811;
		343	:fraction <= 6828;
		344	:fraction <= 6846;
		345	:fraction <= 6863;
		346	:fraction <= 6880;
		347	:fraction <= 6897;
		348	:fraction <= 6915;
		349	:fraction <= 6932;
		350	:fraction <= 6949;
		351	:fraction <= 6966;
		352	:fraction <= 6983;
		353	:fraction <= 7001;
		354	:fraction <= 7018;
		355	:fraction <= 7035;
		356	:fraction <= 7052;
		357	:fraction <= 7069;
		358	:fraction <= 7086;
		359	:fraction <= 7103;
		360	:fraction <= 7120;
		361	:fraction <= 7138;
		362	:fraction <= 7155;
		363	:fraction <= 7172;
		364	:fraction <= 7189;
		365	:fraction <= 7206;
		366	:fraction <= 7223;
		367	:fraction <= 7240;
		368	:fraction <= 7257;
		369	:fraction <= 7274;
		370	:fraction <= 7291;
		371	:fraction <= 7308;
		372	:fraction <= 7325;
		373	:fraction <= 7341;
		374	:fraction <= 7358;
		375	:fraction <= 7375;
		376	:fraction <= 7392;
		377	:fraction <= 7409;
		378	:fraction <= 7426;
		379	:fraction <= 7443;
		380	:fraction <= 7460;
		381	:fraction <= 7476;
		382	:fraction <= 7493;
		383	:fraction <= 7510;
		384	:fraction <= 7527;
		385	:fraction <= 7544;
		386	:fraction <= 7560;
		387	:fraction <= 7577;
		388	:fraction <= 7594;
		389	:fraction <= 7611;
		390	:fraction <= 7627;
		391	:fraction <= 7644;
		392	:fraction <= 7661;
		393	:fraction <= 7677;
		394	:fraction <= 7694;
		395	:fraction <= 7711;
		396	:fraction <= 7727;
		397	:fraction <= 7744;
		398	:fraction <= 7761;
		399	:fraction <= 7777;
		400	:fraction <= 7794;
		401	:fraction <= 7811;
		402	:fraction <= 7827;
		403	:fraction <= 7844;
		404	:fraction <= 7860;
		405	:fraction <= 7877;
		406	:fraction <= 7893;
		407	:fraction <= 7910;
		408	:fraction <= 7926;
		409	:fraction <= 7943;
		410	:fraction <= 7959;
		411	:fraction <= 7976;
		412	:fraction <= 7992;
		413	:fraction <= 8009;
		414	:fraction <= 8025;
		415	:fraction <= 8042;
		416	:fraction <= 8058;
		417	:fraction <= 8074;
		418	:fraction <= 8091;
		419	:fraction <= 8107;
		420	:fraction <= 8124;
		421	:fraction <= 8140;
		422	:fraction <= 8156;
		423	:fraction <= 8173;
		424	:fraction <= 8189;
		425	:fraction <= 8205;
		426	:fraction <= 8222;
		427	:fraction <= 8238;
		428	:fraction <= 8254;
		429	:fraction <= 8270;
		430	:fraction <= 8287;
		431	:fraction <= 8303;
		432	:fraction <= 8319;
		433	:fraction <= 8335;
		434	:fraction <= 8352;
		435	:fraction <= 8368;
		436	:fraction <= 8384;
		437	:fraction <= 8400;
		438	:fraction <= 8416;
		439	:fraction <= 8433;
		440	:fraction <= 8449;
		441	:fraction <= 8465;
		442	:fraction <= 8481;
		443	:fraction <= 8497;
		444	:fraction <= 8513;
		445	:fraction <= 8529;
		446	:fraction <= 8545;
		447	:fraction <= 8561;
		448	:fraction <= 8578;
		449	:fraction <= 8594;
		450	:fraction <= 8610;
		451	:fraction <= 8626;
		452	:fraction <= 8642;
		453	:fraction <= 8658;
		454	:fraction <= 8674;
		455	:fraction <= 8690;
		456	:fraction <= 8706;
		457	:fraction <= 8722;
		458	:fraction <= 8738;
		459	:fraction <= 8754;
		460	:fraction <= 8769;
		461	:fraction <= 8785;
		462	:fraction <= 8801;
		463	:fraction <= 8817;
		464	:fraction <= 8833;
		465	:fraction <= 8849;
		466	:fraction <= 8865;
		467	:fraction <= 8881;
		468	:fraction <= 8897;
		469	:fraction <= 8912;
		470	:fraction <= 8928;
		471	:fraction <= 8944;
		472	:fraction <= 8960;
		473	:fraction <= 8976;
		474	:fraction <= 8991;
		475	:fraction <= 9007;
		476	:fraction <= 9023;
		477	:fraction <= 9039;
		478	:fraction <= 9054;
		479	:fraction <= 9070;
		480	:fraction <= 9086;
		481	:fraction <= 9102;
		482	:fraction <= 9117;
		483	:fraction <= 9133;
		484	:fraction <= 9149;
		485	:fraction <= 9164;
		486	:fraction <= 9180;
		487	:fraction <= 9196;
		488	:fraction <= 9211;
		489	:fraction <= 9227;
		490	:fraction <= 9243;
		491	:fraction <= 9258;
		492	:fraction <= 9274;
		493	:fraction <= 9289;
		494	:fraction <= 9305;
		495	:fraction <= 9320;
		496	:fraction <= 9336;
		497	:fraction <= 9352;
		498	:fraction <= 9367;
		499	:fraction <= 9383;
		500	:fraction <= 9398;
		501	:fraction <= 9414;
		502	:fraction <= 9429;
		503	:fraction <= 9445;
		504	:fraction <= 9460;
		505	:fraction <= 9476;
		506	:fraction <= 9491;
		507	:fraction <= 9506;
		508	:fraction <= 9522;
		509	:fraction <= 9537;
		510	:fraction <= 9553;
		511	:fraction <= 9568;
		512	:fraction <= 9584;
		513	:fraction <= 9599;
		514	:fraction <= 9614;
		515	:fraction <= 9630;
		516	:fraction <= 9645;
		517	:fraction <= 9660;
		518	:fraction <= 9676;
		519	:fraction <= 9691;
		520	:fraction <= 9706;
		521	:fraction <= 9722;
		522	:fraction <= 9737;
		523	:fraction <= 9752;
		524	:fraction <= 9767;
		525	:fraction <= 9783;
		526	:fraction <= 9798;
		527	:fraction <= 9813;
		528	:fraction <= 9828;
		529	:fraction <= 9844;
		530	:fraction <= 9859;
		531	:fraction <= 9874;
		532	:fraction <= 9889;
		533	:fraction <= 9905;
		534	:fraction <= 9920;
		535	:fraction <= 9935;
		536	:fraction <= 9950;
		537	:fraction <= 9965;
		538	:fraction <= 9980;
		539	:fraction <= 9995;
		540	:fraction <= 10011;
		541	:fraction <= 10026;
		542	:fraction <= 10041;
		543	:fraction <= 10056;
		544	:fraction <= 10071;
		545	:fraction <= 10086;
		546	:fraction <= 10101;
		547	:fraction <= 10116;
		548	:fraction <= 10131;
		549	:fraction <= 10146;
		550	:fraction <= 10161;
		551	:fraction <= 10176;
		552	:fraction <= 10191;
		553	:fraction <= 10206;
		554	:fraction <= 10221;
		555	:fraction <= 10236;
		556	:fraction <= 10251;
		557	:fraction <= 10266;
		558	:fraction <= 10281;
		559	:fraction <= 10296;
		560	:fraction <= 10311;
		561	:fraction <= 10326;
		562	:fraction <= 10341;
		563	:fraction <= 10356;
		564	:fraction <= 10370;
		565	:fraction <= 10385;
		566	:fraction <= 10400;
		567	:fraction <= 10415;
		568	:fraction <= 10430;
		569	:fraction <= 10445;
		570	:fraction <= 10460;
		571	:fraction <= 10474;
		572	:fraction <= 10489;
		573	:fraction <= 10504;
		574	:fraction <= 10519;
		575	:fraction <= 10534;
		576	:fraction <= 10548;
		577	:fraction <= 10563;
		578	:fraction <= 10578;
		579	:fraction <= 10593;
		580	:fraction <= 10607;
		581	:fraction <= 10622;
		582	:fraction <= 10637;
		583	:fraction <= 10652;
		584	:fraction <= 10666;
		585	:fraction <= 10681;
		586	:fraction <= 10696;
		587	:fraction <= 10710;
		588	:fraction <= 10725;
		589	:fraction <= 10740;
		590	:fraction <= 10754;
		591	:fraction <= 10769;
		592	:fraction <= 10784;
		593	:fraction <= 10798;
		594	:fraction <= 10813;
		595	:fraction <= 10827;
		596	:fraction <= 10842;
		597	:fraction <= 10857;
		598	:fraction <= 10871;
		599	:fraction <= 10886;
		600	:fraction <= 10900;
		601	:fraction <= 10915;
		602	:fraction <= 10929;
		603	:fraction <= 10944;
		604	:fraction <= 10959;
		605	:fraction <= 10973;
		606	:fraction <= 10988;
		607	:fraction <= 11002;
		608	:fraction <= 11017;
		609	:fraction <= 11031;
		610	:fraction <= 11045;
		611	:fraction <= 11060;
		612	:fraction <= 11074;
		613	:fraction <= 11089;
		614	:fraction <= 11103;
		615	:fraction <= 11118;
		616	:fraction <= 11132;
		617	:fraction <= 11147;
		618	:fraction <= 11161;
		619	:fraction <= 11175;
		620	:fraction <= 11190;
		621	:fraction <= 11204;
		622	:fraction <= 11218;
		623	:fraction <= 11233;
		624	:fraction <= 11247;
		625	:fraction <= 11261;
		626	:fraction <= 11276;
		627	:fraction <= 11290;
		628	:fraction <= 11304;
		629	:fraction <= 11319;
		630	:fraction <= 11333;
		631	:fraction <= 11347;
		632	:fraction <= 11362;
		633	:fraction <= 11376;
		634	:fraction <= 11390;
		635	:fraction <= 11404;
		636	:fraction <= 11419;
		637	:fraction <= 11433;
		638	:fraction <= 11447;
		639	:fraction <= 11461;
		640	:fraction <= 11476;
		641	:fraction <= 11490;
		642	:fraction <= 11504;
		643	:fraction <= 11518;
		644	:fraction <= 11532;
		645	:fraction <= 11546;
		646	:fraction <= 11561;
		647	:fraction <= 11575;
		648	:fraction <= 11589;
		649	:fraction <= 11603;
		650	:fraction <= 11617;
		651	:fraction <= 11631;
		652	:fraction <= 11645;
		653	:fraction <= 11659;
		654	:fraction <= 11674;
		655	:fraction <= 11688;
		656	:fraction <= 11702;
		657	:fraction <= 11716;
		658	:fraction <= 11730;
		659	:fraction <= 11744;
		660	:fraction <= 11758;
		661	:fraction <= 11772;
		662	:fraction <= 11786;
		663	:fraction <= 11800;
		664	:fraction <= 11814;
		665	:fraction <= 11828;
		666	:fraction <= 11842;
		667	:fraction <= 11856;
		668	:fraction <= 11870;
		669	:fraction <= 11884;
		670	:fraction <= 11898;
		671	:fraction <= 11912;
		672	:fraction <= 11926;
		673	:fraction <= 11940;
		674	:fraction <= 11954;
		675	:fraction <= 11968;
		676	:fraction <= 11981;
		677	:fraction <= 11995;
		678	:fraction <= 12009;
		679	:fraction <= 12023;
		680	:fraction <= 12037;
		681	:fraction <= 12051;
		682	:fraction <= 12065;
		683	:fraction <= 12079;
		684	:fraction <= 12092;
		685	:fraction <= 12106;
		686	:fraction <= 12120;
		687	:fraction <= 12134;
		688	:fraction <= 12148;
		689	:fraction <= 12161;
		690	:fraction <= 12175;
		691	:fraction <= 12189;
		692	:fraction <= 12203;
		693	:fraction <= 12217;
		694	:fraction <= 12230;
		695	:fraction <= 12244;
		696	:fraction <= 12258;
		697	:fraction <= 12272;
		698	:fraction <= 12285;
		699	:fraction <= 12299;
		700	:fraction <= 12313;
		701	:fraction <= 12327;
		702	:fraction <= 12340;
		703	:fraction <= 12354;
		704	:fraction <= 12368;
		705	:fraction <= 12381;
		706	:fraction <= 12395;
		707	:fraction <= 12409;
		708	:fraction <= 12422;
		709	:fraction <= 12436;
		710	:fraction <= 12450;
		711	:fraction <= 12463;
		712	:fraction <= 12477;
		713	:fraction <= 12490;
		714	:fraction <= 12504;
		715	:fraction <= 12518;
		716	:fraction <= 12531;
		717	:fraction <= 12545;
		718	:fraction <= 12558;
		719	:fraction <= 12572;
		720	:fraction <= 12585;
		721	:fraction <= 12599;
		722	:fraction <= 12613;
		723	:fraction <= 12626;
		724	:fraction <= 12640;
		725	:fraction <= 12653;
		726	:fraction <= 12667;
		727	:fraction <= 12680;
		728	:fraction <= 12694;
		729	:fraction <= 12707;
		730	:fraction <= 12721;
		731	:fraction <= 12734;
		732	:fraction <= 12748;
		733	:fraction <= 12761;
		734	:fraction <= 12774;
		735	:fraction <= 12788;
		736	:fraction <= 12801;
		737	:fraction <= 12815;
		738	:fraction <= 12828;
		739	:fraction <= 12842;
		740	:fraction <= 12855;
		741	:fraction <= 12868;
		742	:fraction <= 12882;
		743	:fraction <= 12895;
		744	:fraction <= 12908;
		745	:fraction <= 12922;
		746	:fraction <= 12935;
		747	:fraction <= 12949;
		748	:fraction <= 12962;
		749	:fraction <= 12975;
		750	:fraction <= 12989;
		751	:fraction <= 13002;
		752	:fraction <= 13015;
		753	:fraction <= 13029;
		754	:fraction <= 13042;
		755	:fraction <= 13055;
		756	:fraction <= 13068;
		757	:fraction <= 13082;
		758	:fraction <= 13095;
		759	:fraction <= 13108;
		760	:fraction <= 13121;
		761	:fraction <= 13135;
		762	:fraction <= 13148;
		763	:fraction <= 13161;
		764	:fraction <= 13174;
		765	:fraction <= 13188;
		766	:fraction <= 13201;
		767	:fraction <= 13214;
		768	:fraction <= 13227;
		769	:fraction <= 13240;
		770	:fraction <= 13254;
		771	:fraction <= 13267;
		772	:fraction <= 13280;
		773	:fraction <= 13293;
		774	:fraction <= 13306;
		775	:fraction <= 13319;
		776	:fraction <= 13332;
		777	:fraction <= 13346;
		778	:fraction <= 13359;
		779	:fraction <= 13372;
		780	:fraction <= 13385;
		781	:fraction <= 13398;
		782	:fraction <= 13411;
		783	:fraction <= 13424;
		784	:fraction <= 13437;
		785	:fraction <= 13450;
		786	:fraction <= 13463;
		787	:fraction <= 13477;
		788	:fraction <= 13490;
		789	:fraction <= 13503;
		790	:fraction <= 13516;
		791	:fraction <= 13529;
		792	:fraction <= 13542;
		793	:fraction <= 13555;
		794	:fraction <= 13568;
		795	:fraction <= 13581;
		796	:fraction <= 13594;
		797	:fraction <= 13607;
		798	:fraction <= 13620;
		799	:fraction <= 13633;
		800	:fraction <= 13646;
		801	:fraction <= 13659;
		802	:fraction <= 13671;
		803	:fraction <= 13684;
		804	:fraction <= 13697;
		805	:fraction <= 13710;
		806	:fraction <= 13723;
		807	:fraction <= 13736;
		808	:fraction <= 13749;
		809	:fraction <= 13762;
		810	:fraction <= 13775;
		811	:fraction <= 13788;
		812	:fraction <= 13801;
		813	:fraction <= 13813;
		814	:fraction <= 13826;
		815	:fraction <= 13839;
		816	:fraction <= 13852;
		817	:fraction <= 13865;
		818	:fraction <= 13878;
		819	:fraction <= 13891;
		820	:fraction <= 13903;
		821	:fraction <= 13916;
		822	:fraction <= 13929;
		823	:fraction <= 13942;
		824	:fraction <= 13955;
		825	:fraction <= 13967;
		826	:fraction <= 13980;
		827	:fraction <= 13993;
		828	:fraction <= 14006;
		829	:fraction <= 14018;
		830	:fraction <= 14031;
		831	:fraction <= 14044;
		832	:fraction <= 14057;
		833	:fraction <= 14069;
		834	:fraction <= 14082;
		835	:fraction <= 14095;
		836	:fraction <= 14108;
		837	:fraction <= 14120;
		838	:fraction <= 14133;
		839	:fraction <= 14146;
		840	:fraction <= 14158;
		841	:fraction <= 14171;
		842	:fraction <= 14184;
		843	:fraction <= 14196;
		844	:fraction <= 14209;
		845	:fraction <= 14222;
		846	:fraction <= 14234;
		847	:fraction <= 14247;
		848	:fraction <= 14260;
		849	:fraction <= 14272;
		850	:fraction <= 14285;
		851	:fraction <= 14297;
		852	:fraction <= 14310;
		853	:fraction <= 14323;
		854	:fraction <= 14335;
		855	:fraction <= 14348;
		856	:fraction <= 14360;
		857	:fraction <= 14373;
		858	:fraction <= 14385;
		859	:fraction <= 14398;
		860	:fraction <= 14411;
		861	:fraction <= 14423;
		862	:fraction <= 14436;
		863	:fraction <= 14448;
		864	:fraction <= 14461;
		865	:fraction <= 14473;
		866	:fraction <= 14486;
		867	:fraction <= 14498;
		868	:fraction <= 14511;
		869	:fraction <= 14523;
		870	:fraction <= 14536;
		871	:fraction <= 14548;
		872	:fraction <= 14561;
		873	:fraction <= 14573;
		874	:fraction <= 14586;
		875	:fraction <= 14598;
		876	:fraction <= 14610;
		877	:fraction <= 14623;
		878	:fraction <= 14635;
		879	:fraction <= 14648;
		880	:fraction <= 14660;
		881	:fraction <= 14673;
		882	:fraction <= 14685;
		883	:fraction <= 14697;
		884	:fraction <= 14710;
		885	:fraction <= 14722;
		886	:fraction <= 14735;
		887	:fraction <= 14747;
		888	:fraction <= 14759;
		889	:fraction <= 14772;
		890	:fraction <= 14784;
		891	:fraction <= 14796;
		892	:fraction <= 14809;
		893	:fraction <= 14821;
		894	:fraction <= 14833;
		895	:fraction <= 14846;
		896	:fraction <= 14858;
		897	:fraction <= 14870;
		898	:fraction <= 14883;
		899	:fraction <= 14895;
		900	:fraction <= 14907;
		901	:fraction <= 14919;
		902	:fraction <= 14932;
		903	:fraction <= 14944;
		904	:fraction <= 14956;
		905	:fraction <= 14969;
		906	:fraction <= 14981;
		907	:fraction <= 14993;
		908	:fraction <= 15005;
		909	:fraction <= 15017;
		910	:fraction <= 15030;
		911	:fraction <= 15042;
		912	:fraction <= 15054;
		913	:fraction <= 15066;
		914	:fraction <= 15079;
		915	:fraction <= 15091;
		916	:fraction <= 15103;
		917	:fraction <= 15115;
		918	:fraction <= 15127;
		919	:fraction <= 15139;
		920	:fraction <= 15152;
		921	:fraction <= 15164;
		922	:fraction <= 15176;
		923	:fraction <= 15188;
		924	:fraction <= 15200;
		925	:fraction <= 15212;
		926	:fraction <= 15224;
		927	:fraction <= 15237;
		928	:fraction <= 15249;
		929	:fraction <= 15261;
		930	:fraction <= 15273;
		931	:fraction <= 15285;
		932	:fraction <= 15297;
		933	:fraction <= 15309;
		934	:fraction <= 15321;
		935	:fraction <= 15333;
		936	:fraction <= 15345;
		937	:fraction <= 15357;
		938	:fraction <= 15369;
		939	:fraction <= 15382;
		940	:fraction <= 15394;
		941	:fraction <= 15406;
		942	:fraction <= 15418;
		943	:fraction <= 15430;
		944	:fraction <= 15442;
		945	:fraction <= 15454;
		946	:fraction <= 15466;
		947	:fraction <= 15478;
		948	:fraction <= 15490;
		949	:fraction <= 15502;
		950	:fraction <= 15514;
		951	:fraction <= 15526;
		952	:fraction <= 15538;
		953	:fraction <= 15550;
		954	:fraction <= 15561;
		955	:fraction <= 15573;
		956	:fraction <= 15585;
		957	:fraction <= 15597;
		958	:fraction <= 15609;
		959	:fraction <= 15621;
		960	:fraction <= 15633;
		961	:fraction <= 15645;
		962	:fraction <= 15657;
		963	:fraction <= 15669;
		964	:fraction <= 15681;
		965	:fraction <= 15693;
		966	:fraction <= 15704;
		967	:fraction <= 15716;
		968	:fraction <= 15728;
		969	:fraction <= 15740;
		970	:fraction <= 15752;
		971	:fraction <= 15764;
		972	:fraction <= 15776;
		973	:fraction <= 15787;
		974	:fraction <= 15799;
		975	:fraction <= 15811;
		976	:fraction <= 15823;
		977	:fraction <= 15835;
		978	:fraction <= 15847;
		979	:fraction <= 15858;
		980	:fraction <= 15870;
		981	:fraction <= 15882;
		982	:fraction <= 15894;
		983	:fraction <= 15905;
		984	:fraction <= 15917;
		985	:fraction <= 15929;
		986	:fraction <= 15941;
		987	:fraction <= 15953;
		988	:fraction <= 15964;
		989	:fraction <= 15976;
		990	:fraction <= 15988;
		991	:fraction <= 16000;
		992	:fraction <= 16011;
		993	:fraction <= 16023;
		994	:fraction <= 16035;
		995	:fraction <= 16046;
		996	:fraction <= 16058;
		997	:fraction <= 16070;
		998	:fraction <= 16081;
		999	:fraction <= 16093;
		1000	:fraction <= 16105;
		1001	:fraction <= 16117;
		1002	:fraction <= 16128;
		1003	:fraction <= 16140;
		1004	:fraction <= 16152;
		1005	:fraction <= 16163;
		1006	:fraction <= 16175;
		1007	:fraction <= 16186;
		1008	:fraction <= 16198;
		1009	:fraction <= 16210;
		1010	:fraction <= 16221;
		1011	:fraction <= 16233;
		1012	:fraction <= 16245;
		1013	:fraction <= 16256;
		1014	:fraction <= 16268;
		1015	:fraction <= 16279;
		1016	:fraction <= 16291;
		1017	:fraction <= 16303;
		1018	:fraction <= 16314;
		1019	:fraction <= 16326;
		1020	:fraction <= 16337;
		1021	:fraction <= 16349;
		1022	:fraction <= 16360;
		1023	:fraction <= 16372;
		 endcase
	      end
	      4:begin
		 //! Output Data
		 outdata<=inte*16384+fraction;
		 dv<=1;
	      end
	    endcase

	 end // else: !if(inte==0)
      end else begin // if (start==1)
	 /* Offline  */
	 clk_cnt<=0;
	 dv<=0;
	 inte<=63;
      end // else: !if(start==1)
   end // always@ (posedge clk)
   

endmodule
